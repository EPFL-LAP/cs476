module biosRom ( input wire        clock,
                 input wire [11:0] address,
                 output reg [31:0] romData);

  always @*
    case (address)
      12'b000000000000 : romData <= 32'h0013ADDE;
      12'b000000000001 : romData <= 32'h00000015;
      12'b000000000010 : romData <= 32'h21000000;
      12'b000000000011 : romData <= 32'h00000015;
      12'b000000000100 : romData <= 32'h1F000000;
      12'b000000000101 : romData <= 32'h00000015;
      12'b000000000110 : romData <= 32'h1D000000;
      12'b000000000111 : romData <= 32'h00000015;
      12'b000000001000 : romData <= 32'h1B000000;
      12'b000000001001 : romData <= 32'h00000015;
      12'b000000001010 : romData <= 32'h19000000;
      12'b000000001011 : romData <= 32'h00000015;
      12'b000000001100 : romData <= 32'h17000000;
      12'b000000001101 : romData <= 32'h00000015;
      12'b000000001110 : romData <= 32'h15000000;
      12'b000000001111 : romData <= 32'h00000015;
      12'b000000010000 : romData <= 32'h13000000;
      12'b000000010001 : romData <= 32'h00000015;
      12'b000000010010 : romData <= 32'h11000000;
      12'b000000010011 : romData <= 32'h00000015;
      12'b000000010100 : romData <= 32'h0F000000;
      12'b000000010101 : romData <= 32'h00000015;
      12'b000000010110 : romData <= 32'h0D000000;
      12'b000000010111 : romData <= 32'h00000015;
      12'b000000011000 : romData <= 32'h0B000000;
      12'b000000011001 : romData <= 32'h00000015;
      12'b000000011010 : romData <= 32'h09000000;
      12'b000000011011 : romData <= 32'h00000015;
      12'b000000011100 : romData <= 32'h00C02018;
      12'b000000011101 : romData <= 32'hFC1F21A8;
      12'b000000011110 : romData <= 32'h050060E0;
      12'b000000011111 : romData <= 32'hE4030004;
      12'b000000100000 : romData <= 32'h050080E0;
      12'b000000100010 : romData <= 32'h00000015;
      12'b000000100011 : romData <= 32'h84FF219C;
      12'b000000100100 : romData <= 32'h001001D4;
      12'b000000100101 : romData <= 32'h041801D4;
      12'b000000100110 : romData <= 32'h082001D4;
      12'b000000100111 : romData <= 32'h0C2801D4;
      12'b000000101000 : romData <= 32'h103001D4;
      12'b000000101001 : romData <= 32'h143801D4;
      12'b000000101010 : romData <= 32'h184001D4;
      12'b000000101011 : romData <= 32'h1C4801D4;
      12'b000000101100 : romData <= 32'h205001D4;
      12'b000000101101 : romData <= 32'h245801D4;
      12'b000000101110 : romData <= 32'h286001D4;
      12'b000000101111 : romData <= 32'h2C6801D4;
      12'b000000110000 : romData <= 32'h307001D4;
      12'b000000110001 : romData <= 32'h347801D4;
      12'b000000110010 : romData <= 32'h388001D4;
      12'b000000110011 : romData <= 32'h3C8801D4;
      12'b000000110100 : romData <= 32'h409001D4;
      12'b000000110101 : romData <= 32'h449801D4;
      12'b000000110110 : romData <= 32'h48A001D4;
      12'b000000110111 : romData <= 32'h4CA801D4;
      12'b000000111000 : romData <= 32'h50B001D4;
      12'b000000111001 : romData <= 32'h54B801D4;
      12'b000000111010 : romData <= 32'h58C001D4;
      12'b000000111011 : romData <= 32'h5CC801D4;
      12'b000000111100 : romData <= 32'h60D001D4;
      12'b000000111101 : romData <= 32'h64D801D4;
      12'b000000111110 : romData <= 32'h68E001D4;
      12'b000000111111 : romData <= 32'h6CE801D4;
      12'b000001000000 : romData <= 32'h70F001D4;
      12'b000001000001 : romData <= 32'h74F801D4;
      12'b000001000010 : romData <= 32'h1200E0B7;
      12'b000001000011 : romData <= 32'h0200FFBB;
      12'b000001000100 : romData <= 32'h00F0C01B;
      12'b000001000101 : romData <= 32'hAC01DEAB;
      12'b000001000110 : romData <= 32'h00F8DEE3;
      12'b000001000111 : romData <= 32'h0000FE87;
      12'b000001001000 : romData <= 32'h00F80048;
      12'b000001001001 : romData <= 32'h00000015;
      12'b000001001010 : romData <= 32'h00004184;
      12'b000001001011 : romData <= 32'h04006184;
      12'b000001001100 : romData <= 32'h08008184;
      12'b000001001101 : romData <= 32'h0C00A184;
      12'b000001001110 : romData <= 32'h1000C184;
      12'b000001001111 : romData <= 32'h1400E184;
      12'b000001010000 : romData <= 32'h18000185;
      12'b000001010001 : romData <= 32'h1C002185;
      12'b000001010010 : romData <= 32'h20004185;
      12'b000001010011 : romData <= 32'h24006185;
      12'b000001010100 : romData <= 32'h28008185;
      12'b000001010101 : romData <= 32'h2C00A185;
      12'b000001010110 : romData <= 32'h3000C185;
      12'b000001010111 : romData <= 32'h3400E185;
      12'b000001011000 : romData <= 32'h38000186;
      12'b000001011001 : romData <= 32'h3C002186;
      12'b000001011010 : romData <= 32'h40004186;
      12'b000001011011 : romData <= 32'h44006186;
      12'b000001011100 : romData <= 32'h48008186;
      12'b000001011101 : romData <= 32'h4C00A186;
      12'b000001011110 : romData <= 32'h5000C186;
      12'b000001011111 : romData <= 32'h5400E186;
      12'b000001100000 : romData <= 32'h58000187;
      12'b000001100001 : romData <= 32'h5C002187;
      12'b000001100010 : romData <= 32'h60004187;
      12'b000001100011 : romData <= 32'h64006187;
      12'b000001100100 : romData <= 32'h68008187;
      12'b000001100101 : romData <= 32'h6C00A187;
      12'b000001100110 : romData <= 32'h7000C187;
      12'b000001100111 : romData <= 32'h7400E187;
      12'b000001101000 : romData <= 32'h7C00219C;
      12'b000001101001 : romData <= 32'h00000024;
      12'b000001101010 : romData <= 32'h00000015;
      12'b000001101011 : romData <= 32'h700000F0;
      12'b000001101100 : romData <= 32'hE40100F0;
      12'b000001101101 : romData <= 32'h000200F0;
      12'b000001101110 : romData <= 32'h1C0200F0;
      12'b000001101111 : romData <= 32'h380200F0;
      12'b000001110000 : romData <= 32'h540200F0;
      12'b000001110001 : romData <= 32'h700200F0;
      12'b000001110010 : romData <= 32'h8C0200F0;
      12'b000001110011 : romData <= 32'hA80200F0;
      12'b000001110100 : romData <= 32'hC40200F0;
      12'b000001110101 : romData <= 32'hE00200F0;
      12'b000001110110 : romData <= 32'hFC0200F0;
      12'b000001110111 : romData <= 32'h340300F0;
      12'b000001111000 : romData <= 32'h180300F0;
      12'b000001111001 : romData <= 32'h00F0A018;
      12'b000001111010 : romData <= 32'h00F08018;
      12'b000001111011 : romData <= 32'h00F06018;
      12'b000001111100 : romData <= 32'hF01CA59C;
      12'b000001111101 : romData <= 32'h7809849C;
      12'b000001111110 : romData <= 32'h5D010000;
      12'b000001111111 : romData <= 32'hD00A639C;
      12'b000010000000 : romData <= 32'h00F0A018;
      12'b000010000001 : romData <= 32'h00F08018;
      12'b000010000010 : romData <= 32'h00F06018;
      12'b000010000011 : romData <= 32'hFC1CA59C;
      12'b000010000100 : romData <= 32'h7809849C;
      12'b000010000101 : romData <= 32'h56010000;
      12'b000010000110 : romData <= 32'hD00A639C;
      12'b000010000111 : romData <= 32'h00F0A018;
      12'b000010001000 : romData <= 32'h00F08018;
      12'b000010001001 : romData <= 32'h00F06018;
      12'b000010001010 : romData <= 32'h0D1DA59C;
      12'b000010001011 : romData <= 32'h7809849C;
      12'b000010001100 : romData <= 32'h4F010000;
      12'b000010001101 : romData <= 32'hD00A639C;
      12'b000010001110 : romData <= 32'h00F0A018;
      12'b000010001111 : romData <= 32'h00F08018;
      12'b000010010000 : romData <= 32'h00F06018;
      12'b000010010001 : romData <= 32'h1B1DA59C;
      12'b000010010010 : romData <= 32'h7809849C;
      12'b000010010011 : romData <= 32'h48010000;
      12'b000010010100 : romData <= 32'hD00A639C;
      12'b000010010101 : romData <= 32'h00F0A018;
      12'b000010010110 : romData <= 32'h00F08018;
      12'b000010010111 : romData <= 32'h00F06018;
      12'b000010011000 : romData <= 32'h211DA59C;
      12'b000010011001 : romData <= 32'h7809849C;
      12'b000010011010 : romData <= 32'h41010000;
      12'b000010011011 : romData <= 32'hD00A639C;
      12'b000010011100 : romData <= 32'h00F0A018;
      12'b000010011101 : romData <= 32'h00F08018;
      12'b000010011110 : romData <= 32'h00F06018;
      12'b000010011111 : romData <= 32'h2A1DA59C;
      12'b000010100000 : romData <= 32'h7809849C;
      12'b000010100001 : romData <= 32'h3A010000;
      12'b000010100010 : romData <= 32'hD00A639C;
      12'b000010100011 : romData <= 32'h00F0A018;
      12'b000010100100 : romData <= 32'h00F08018;
      12'b000010100101 : romData <= 32'h00F06018;
      12'b000010100110 : romData <= 32'h301DA59C;
      12'b000010100111 : romData <= 32'h7809849C;
      12'b000010101000 : romData <= 32'h33010000;
      12'b000010101001 : romData <= 32'hD00A639C;
      12'b000010101010 : romData <= 32'h00F0A018;
      12'b000010101011 : romData <= 32'h00F08018;
      12'b000010101100 : romData <= 32'h00F06018;
      12'b000010101101 : romData <= 32'h361DA59C;
      12'b000010101110 : romData <= 32'h7809849C;
      12'b000010101111 : romData <= 32'h2C010000;
      12'b000010110000 : romData <= 32'hD00A639C;
      12'b000010110001 : romData <= 32'h00F0A018;
      12'b000010110010 : romData <= 32'h00F08018;
      12'b000010110011 : romData <= 32'h00F06018;
      12'b000010110100 : romData <= 32'h3C1DA59C;
      12'b000010110101 : romData <= 32'h7809849C;
      12'b000010110110 : romData <= 32'h25010000;
      12'b000010110111 : romData <= 32'hD00A639C;
      12'b000010111000 : romData <= 32'h00F0A018;
      12'b000010111001 : romData <= 32'h00F08018;
      12'b000010111010 : romData <= 32'h00F06018;
      12'b000010111011 : romData <= 32'h421DA59C;
      12'b000010111100 : romData <= 32'h7809849C;
      12'b000010111101 : romData <= 32'h1E010000;
      12'b000010111110 : romData <= 32'hD00A639C;
      12'b000010111111 : romData <= 32'h00F0A018;
      12'b000011000000 : romData <= 32'h00F08018;
      12'b000011000001 : romData <= 32'h00F06018;
      12'b000011000010 : romData <= 32'h4A1DA59C;
      12'b000011000011 : romData <= 32'h7809849C;
      12'b000011000100 : romData <= 32'h17010000;
      12'b000011000101 : romData <= 32'hD00A639C;
      12'b000011000110 : romData <= 32'h00F0A018;
      12'b000011000111 : romData <= 32'h00F08018;
      12'b000011001000 : romData <= 32'h00F06018;
      12'b000011001001 : romData <= 32'h531DA59C;
      12'b000011001010 : romData <= 32'h7809849C;
      12'b000011001011 : romData <= 32'h10010000;
      12'b000011001100 : romData <= 32'hD00A639C;
      12'b000011001101 : romData <= 32'h00F0A018;
      12'b000011001110 : romData <= 32'h00F08018;
      12'b000011001111 : romData <= 32'h00F06018;
      12'b000011010000 : romData <= 32'h5A1DA59C;
      12'b000011010001 : romData <= 32'h7809849C;
      12'b000011010010 : romData <= 32'h09010000;
      12'b000011010011 : romData <= 32'hD00A639C;
      12'b000011010100 : romData <= 32'h0000601A;
      12'b000011010101 : romData <= 32'h0700A0AA;
      12'b000011010110 : romData <= 32'h02A83372;
      12'b000011010111 : romData <= 32'h0000E01A;
      12'b000011011000 : romData <= 32'h010031A6;
      12'b000011011001 : romData <= 32'h00B831E4;
      12'b000011011010 : romData <= 32'hFCFFFF13;
      12'b000011011011 : romData <= 32'h00000015;
      12'b000011011100 : romData <= 32'h00480044;
      12'b000011011101 : romData <= 32'h00000015;
      12'b000011011110 : romData <= 32'h00006019;
      12'b000011011111 : romData <= 32'h02186B71;
      12'b000011100000 : romData <= 32'h00480044;
      12'b000011100001 : romData <= 32'h00000015;
      12'b000011100010 : romData <= 32'h160020AA;
      12'b000011100011 : romData <= 32'h02890370;
      12'b000011100100 : romData <= 32'h020020AA;
      12'b000011100101 : romData <= 32'h070060AA;
      12'b000011100110 : romData <= 32'h02991170;
      12'b000011100111 : romData <= 32'hEDFFFF03;
      12'b000011101000 : romData <= 32'h00000015;
      12'b000011101001 : romData <= 32'hE0FF219C;
      12'b000011101010 : romData <= 32'h088001D4;
      12'b000011101011 : romData <= 32'h0C9001D4;
      12'b000011101100 : romData <= 32'h10A001D4;
      12'b000011101101 : romData <= 32'h14B001D4;
      12'b000011101110 : romData <= 32'h18C001D4;
      12'b000011101111 : romData <= 32'h1C4801D4;
      12'b000011110000 : romData <= 32'h0000001A;
      12'b000011110001 : romData <= 32'h0000401A;
      12'b000011110010 : romData <= 32'h160080AA;
      12'b000011110011 : romData <= 32'h0100C0AA;
      12'b000011110100 : romData <= 32'h070000AB;
      12'b000011110101 : romData <= 32'h002092E5;
      12'b000011110110 : romData <= 32'h09000010;
      12'b000011110111 : romData <= 32'h1C002185;
      12'b000011111000 : romData <= 32'h08000186;
      12'b000011111001 : romData <= 32'h0C004186;
      12'b000011111010 : romData <= 32'h10008186;
      12'b000011111011 : romData <= 32'h1400C186;
      12'b000011111100 : romData <= 32'h18000187;
      12'b000011111101 : romData <= 32'h00480044;
      12'b000011111110 : romData <= 32'h2000219C;
      12'b000011111111 : romData <= 32'h02A11070;
      12'b000100000000 : romData <= 32'h180020AA;
      12'b000100000001 : romData <= 32'h008063E2;
      12'b000100000010 : romData <= 32'h0000B386;
      12'b000100000011 : romData <= 32'h0102B572;
      12'b000100000100 : romData <= 32'h02891570;
      12'b000100000101 : romData <= 32'h2000A0AA;
      12'b000100000110 : romData <= 32'h0100319E;
      12'b000100000111 : romData <= 32'h00A831E4;
      12'b000100001000 : romData <= 32'hFAFFFF13;
      12'b000100001001 : romData <= 32'h0400739E;
      12'b000100001010 : romData <= 32'h042001D4;
      12'b000100001011 : romData <= 32'h001801D4;
      12'b000100001100 : romData <= 32'h02C11670;
      12'b000100001101 : romData <= 32'hC7FFFF07;
      12'b000100001110 : romData <= 32'h0800529E;
      12'b000100001111 : romData <= 32'h2000109E;
      12'b000100010000 : romData <= 32'h04008184;
      12'b000100010001 : romData <= 32'hE4FFFF03;
      12'b000100010010 : romData <= 32'h00006184;
      12'b000100010011 : romData <= 32'hB8FF219C;
      12'b000100010100 : romData <= 32'h00F08018;
      12'b000100010101 : romData <= 32'h2000A0A8;
      12'b000100010110 : romData <= 32'h8C25849C;
      12'b000100010111 : romData <= 32'h1000619C;
      12'b000100011000 : romData <= 32'h308001D4;
      12'b000100011001 : romData <= 32'h349001D4;
      12'b000100011010 : romData <= 32'h3CB001D4;
      12'b000100011011 : romData <= 32'h40C001D4;
      12'b000100011100 : romData <= 32'h444801D4;
      12'b000100011101 : romData <= 32'h38A001D4;
      12'b000100011110 : romData <= 32'h9B010004;
      12'b000100011111 : romData <= 32'h00F0401A;
      12'b000100100000 : romData <= 32'h00F0001A;
      12'b000100100001 : romData <= 32'h7809529E;
      12'b000100100010 : romData <= 32'hD00A109E;
      12'b000100100011 : romData <= 32'h00F0A018;
      12'b000100100100 : romData <= 32'h611DA59C;
      12'b000100100101 : romData <= 32'h049092E0;
      12'b000100100110 : romData <= 32'hB5000004;
      12'b000100100111 : romData <= 32'h048070E0;
      12'b000100101000 : romData <= 32'h1F00201A;
      12'b000100101001 : romData <= 32'h00F0A018;
      12'b000100101010 : romData <= 32'h0000601A;
      12'b000100101011 : romData <= 32'h00FC31AA;
      12'b000100101100 : romData <= 32'h0004001B;
      12'b000100101101 : romData <= 32'h2000C01A;
      12'b000100101110 : romData <= 32'h921DA59C;
      12'b000100101111 : romData <= 32'h0200A0AA;
      12'b000100110000 : romData <= 32'h08A891E2;
      12'b000100110001 : romData <= 32'h00C094E2;
      12'b000100110010 : romData <= 32'hFFFFE0AE;
      12'b000100110011 : romData <= 32'h0000B486;
      12'b000100110100 : romData <= 32'h00B815E4;
      12'b000100110101 : romData <= 32'h1C000010;
      12'b000100110110 : romData <= 32'h00000015;
      12'b000100110111 : romData <= 32'h0000201A;
      12'b000100111000 : romData <= 32'h008813E4;
      12'b000100111001 : romData <= 32'h0E000010;
      12'b000100111010 : romData <= 32'h049092E0;
      12'b000100111011 : romData <= 32'h00F0A018;
      12'b000100111100 : romData <= 32'h841DA59C;
      12'b000100111101 : romData <= 32'h049092E0;
      12'b000100111110 : romData <= 32'h048070E0;
      12'b000100111111 : romData <= 32'h34004186;
      12'b000101000000 : romData <= 32'h30000186;
      12'b000101000001 : romData <= 32'h38008186;
      12'b000101000010 : romData <= 32'h3C00C186;
      12'b000101000011 : romData <= 32'h40000187;
      12'b000101000100 : romData <= 32'h44002185;
      12'b000101000101 : romData <= 32'h96000000;
      12'b000101000110 : romData <= 32'h4800219C;
      12'b000101000111 : romData <= 32'h048070E0;
      12'b000101001000 : romData <= 32'h93000004;
      12'b000101001001 : romData <= 32'h0C2801D4;
      12'b000101001010 : romData <= 32'h98FFFF07;
      12'b000101001011 : romData <= 32'h04A074E0;
      12'b000101001100 : romData <= 32'h1F00201A;
      12'b000101001101 : romData <= 32'h01FC31AA;
      12'b000101001110 : romData <= 32'h010060AA;
      12'b000101001111 : romData <= 32'hE0FFFF03;
      12'b000101010000 : romData <= 32'h0C00A184;
      12'b000101010001 : romData <= 32'h0100319E;
      12'b000101010010 : romData <= 32'h00B011E4;
      12'b000101010011 : romData <= 32'hDDFFFF0F;
      12'b000101010100 : romData <= 32'h0200A0AA;
      12'b000101010101 : romData <= 32'h00F0A018;
      12'b000101010110 : romData <= 32'hAE1DA59C;
      12'b000101010111 : romData <= 32'h049092E0;
      12'b000101011000 : romData <= 32'h83000004;
      12'b000101011001 : romData <= 32'h048070E0;
      12'b000101011010 : romData <= 32'h1000819E;
      12'b000101011011 : romData <= 32'h04A074E2;
      12'b000101011100 : romData <= 32'h180020AA;
      12'b000101011101 : romData <= 32'h0000B386;
      12'b000101011110 : romData <= 32'h0102B572;
      12'b000101011111 : romData <= 32'h02891570;
      12'b000101100000 : romData <= 32'h2000A0AA;
      12'b000101100001 : romData <= 32'h0100319E;
      12'b000101100010 : romData <= 32'h00A831E4;
      12'b000101100011 : romData <= 32'hFAFFFF13;
      12'b000101100100 : romData <= 32'h0400739E;
      12'b000101100101 : romData <= 32'h7F00201A;
      12'b000101100110 : romData <= 32'h00F031AA;
      12'b000101100111 : romData <= 32'h160060AA;
      12'b000101101000 : romData <= 32'h02991170;
      12'b000101101001 : romData <= 32'h010020AA;
      12'b000101101010 : romData <= 32'h070060AA;
      12'b000101101011 : romData <= 32'h02991170;
      12'b000101101100 : romData <= 32'h68FFFF07;
      12'b000101101101 : romData <= 32'h00000015;
      12'b000101101110 : romData <= 32'h00F0A018;
      12'b000101101111 : romData <= 32'hCF1DA59C;
      12'b000101110000 : romData <= 32'h049092E0;
      12'b000101110001 : romData <= 32'h6A000004;
      12'b000101110010 : romData <= 32'h048070E0;
      12'b000101110011 : romData <= 32'h7F04201A;
      12'b000101110100 : romData <= 32'h00F031AA;
      12'b000101110101 : romData <= 32'h0000601A;
      12'b000101110110 : romData <= 32'h0000B186;
      12'b000101110111 : romData <= 32'h0000F486;
      12'b000101111000 : romData <= 32'h00A817E4;
      12'b000101111001 : romData <= 32'h13000010;
      12'b000101111010 : romData <= 32'h0100739E;
      12'b000101111011 : romData <= 32'hFFFF739E;
      12'b000101111100 : romData <= 32'h00F0A018;
      12'b000101111101 : romData <= 32'h08B801D4;
      12'b000101111110 : romData <= 32'h04A801D4;
      12'b000101111111 : romData <= 32'h009801D4;
      12'b000110000000 : romData <= 32'h049092E0;
      12'b000110000001 : romData <= 32'h048070E0;
      12'b000110000010 : romData <= 32'h59000004;
      12'b000110000011 : romData <= 32'hF41DA59C;
      12'b000110000100 : romData <= 32'h44002185;
      12'b000110000101 : romData <= 32'h30000186;
      12'b000110000110 : romData <= 32'h34004186;
      12'b000110000111 : romData <= 32'h38008186;
      12'b000110001000 : romData <= 32'h3C00C186;
      12'b000110001001 : romData <= 32'h40000187;
      12'b000110001010 : romData <= 32'h00480044;
      12'b000110001011 : romData <= 32'h4800219C;
      12'b000110001100 : romData <= 32'h0800A0AA;
      12'b000110001101 : romData <= 32'h00A833E4;
      12'b000110001110 : romData <= 32'h0400319E;
      12'b000110001111 : romData <= 32'hE7FFFF13;
      12'b000110010000 : romData <= 32'h0400949E;
      12'b000110010001 : romData <= 32'h00F0A018;
      12'b000110010010 : romData <= 32'hABFFFF03;
      12'b000110010011 : romData <= 32'h141EA59C;
      12'b000110010100 : romData <= 32'hF0FF219C;
      12'b000110010101 : romData <= 32'h048001D4;
      12'b000110010110 : romData <= 32'h089001D4;
      12'b000110010111 : romData <= 32'h0C4801D4;
      12'b000110011000 : romData <= 32'h041843E2;
      12'b000110011001 : romData <= 32'h1C0000AA;
      12'b000110011010 : romData <= 32'h488024E2;
      12'b000110011011 : romData <= 32'h0F0031A6;
      12'b000110011100 : romData <= 32'h090060AA;
      12'b000110011101 : romData <= 32'h009851E4;
      12'b000110011110 : romData <= 32'h03000010;
      12'b000110011111 : romData <= 32'h3700719C;
      12'b000110100000 : romData <= 32'h3000719C;
      12'b000110100001 : romData <= 32'h00900048;
      12'b000110100010 : romData <= 32'h002001D4;
      12'b000110100011 : romData <= 32'hFCFF109E;
      12'b000110100100 : romData <= 32'hFCFF20AE;
      12'b000110100101 : romData <= 32'h008830E4;
      12'b000110100110 : romData <= 32'hF4FFFF13;
      12'b000110100111 : romData <= 32'h00008184;
      12'b000110101000 : romData <= 32'h04000186;
      12'b000110101001 : romData <= 32'h08004186;
      12'b000110101010 : romData <= 32'h0C002185;
      12'b000110101011 : romData <= 32'h00480044;
      12'b000110101100 : romData <= 32'h1000219C;
      12'b000110101101 : romData <= 32'hE4FF219C;
      12'b000110101110 : romData <= 32'h0C8001D4;
      12'b000110101111 : romData <= 32'h109001D4;
      12'b000110110000 : romData <= 32'h14A001D4;
      12'b000110110001 : romData <= 32'h184801D4;
      12'b000110110010 : romData <= 32'h041843E2;
      12'b000110110011 : romData <= 32'h0000601A;
      12'b000110110100 : romData <= 32'h0000001A;
      12'b000110110101 : romData <= 32'h0200819E;
      12'b000110110110 : romData <= 32'h0A00A0AA;
      12'b000110110111 : romData <= 32'h0AAB24E3;
      12'b000110111000 : romData <= 32'h020020AA;
      12'b000110111001 : romData <= 32'h088839E2;
      12'b000110111010 : romData <= 32'h00C831E2;
      12'b000110111011 : romData <= 32'h008831E2;
      12'b000110111100 : romData <= 32'h028824E2;
      12'b000110111101 : romData <= 32'h3000319E;
      12'b000110111110 : romData <= 32'h0098F4E2;
      12'b000110111111 : romData <= 32'h008817D8;
      12'b000111000000 : romData <= 32'h0000201A;
      12'b000111000001 : romData <= 32'h008813E4;
      12'b000111000010 : romData <= 32'h04000010;
      12'b000111000011 : romData <= 32'h008804E4;
      12'b000111000100 : romData <= 32'h04000010;
      12'b000111000101 : romData <= 32'h00000015;
      12'b000111000110 : romData <= 32'h0100109E;
      12'b000111000111 : romData <= 32'hFF0010A6;
      12'b000111001000 : romData <= 32'h0100739E;
      12'b000111001001 : romData <= 32'h00A833E4;
      12'b000111001010 : romData <= 32'hEDFFFF13;
      12'b000111001011 : romData <= 32'h0AAB84E0;
      12'b000111001100 : romData <= 32'h0000201A;
      12'b000111001101 : romData <= 32'h008830E4;
      12'b000111001110 : romData <= 32'h07000010;
      12'b000111001111 : romData <= 32'h18002185;
      12'b000111010000 : romData <= 32'h0C000186;
      12'b000111010001 : romData <= 32'h10004186;
      12'b000111010010 : romData <= 32'h14008186;
      12'b000111010011 : romData <= 32'h00480044;
      12'b000111010100 : romData <= 32'h1C00219C;
      12'b000111010101 : romData <= 32'hFFFF109E;
      12'b000111010110 : romData <= 32'h008034E2;
      12'b000111010111 : romData <= 32'h00900048;
      12'b000111011000 : romData <= 32'h0000718C;
      12'b000111011001 : romData <= 32'hF4FFFF03;
      12'b000111011010 : romData <= 32'h0000201A;
      12'b000111011011 : romData <= 32'hE4FF219C;
      12'b000111011100 : romData <= 32'h008001D4;
      12'b000111011101 : romData <= 32'h049001D4;
      12'b000111011110 : romData <= 32'h08A001D4;
      12'b000111011111 : romData <= 32'h0CB001D4;
      12'b000111100000 : romData <= 32'h14D001D4;
      12'b000111100001 : romData <= 32'h10C001D4;
      12'b000111100010 : romData <= 32'h184801D4;
      12'b000111100011 : romData <= 32'h041883E2;
      12'b000111100100 : romData <= 32'h042004E2;
      12'b000111100101 : romData <= 32'h042845E2;
      12'b000111100110 : romData <= 32'h1C00C19E;
      12'b000111100111 : romData <= 32'h250040AB;
      12'b000111101000 : romData <= 32'h00001293;
      12'b000111101001 : romData <= 32'h0000201A;
      12'b000111101010 : romData <= 32'h008838E4;
      12'b000111101011 : romData <= 32'h3C00000C;
      12'b000111101100 : romData <= 32'h00D038E4;
      12'b000111101101 : romData <= 32'h5B000010;
      12'b000111101110 : romData <= 32'h630060AA;
      12'b000111101111 : romData <= 32'h01003292;
      12'b000111110000 : romData <= 32'h009811E4;
      12'b000111110001 : romData <= 32'h4E000010;
      12'b000111110010 : romData <= 32'h009851E5;
      12'b000111110011 : romData <= 32'h1B000010;
      12'b000111110100 : romData <= 32'h0000601A;
      12'b000111110101 : romData <= 32'h009811E4;
      12'b000111110110 : romData <= 32'h29000010;
      12'b000111110111 : romData <= 32'h580060AA;
      12'b000111111000 : romData <= 32'h009811E4;
      12'b000111111001 : romData <= 32'h37000010;
      12'b000111111010 : romData <= 32'h00000015;
      12'b000111111011 : romData <= 32'h00A00048;
      12'b000111111100 : romData <= 32'h250060A8;
      12'b000111111101 : romData <= 32'h0000201A;
      12'b000111111110 : romData <= 32'h008810E4;
      12'b000111111111 : romData <= 32'h04000010;
      12'b001000000000 : romData <= 32'h00000015;
      12'b001000000001 : romData <= 32'h00800048;
      12'b001000000010 : romData <= 32'h250060A8;
      12'b001000000011 : romData <= 32'h0100128F;
      12'b001000000100 : romData <= 32'h00A00048;
      12'b001000000101 : romData <= 32'h04C078E0;
      12'b001000000110 : romData <= 32'h0000201A;
      12'b001000000111 : romData <= 32'h008810E4;
      12'b001000001000 : romData <= 32'h34000010;
      12'b001000001001 : romData <= 32'h00000015;
      12'b001000001010 : romData <= 32'h00800048;
      12'b001000001011 : romData <= 32'h04C078E0;
      12'b001000001100 : romData <= 32'h31000000;
      12'b001000001101 : romData <= 32'h0100529E;
      12'b001000001110 : romData <= 32'h640060AA;
      12'b001000001111 : romData <= 32'h009811E4;
      12'b001000010000 : romData <= 32'hEBFFFF0F;
      12'b001000010001 : romData <= 32'h00000015;
      12'b001000010010 : romData <= 32'h0400169F;
      12'b001000010011 : romData <= 32'h04A074E0;
      12'b001000010100 : romData <= 32'h0000D686;
      12'b001000010101 : romData <= 32'h98FFFF07;
      12'b001000010110 : romData <= 32'h04B096E0;
      12'b001000010111 : romData <= 32'h0000201A;
      12'b001000011000 : romData <= 32'h008810E4;
      12'b001000011001 : romData <= 32'h22000010;
      12'b001000011010 : romData <= 32'h04B096E0;
      12'b001000011011 : romData <= 32'h92FFFF07;
      12'b001000011100 : romData <= 32'h048070E0;
      12'b001000011101 : romData <= 32'h1F000000;
      12'b001000011110 : romData <= 32'h04C0D8E2;
      12'b001000011111 : romData <= 32'h00A00048;
      12'b001000100000 : romData <= 32'h04D07AE0;
      12'b001000100001 : romData <= 32'h0000201A;
      12'b001000100010 : romData <= 32'h008810E4;
      12'b001000100011 : romData <= 32'h04000010;
      12'b001000100100 : romData <= 32'h04D07AE0;
      12'b001000100101 : romData <= 32'h00800048;
      12'b001000100110 : romData <= 32'h00000015;
      12'b001000100111 : romData <= 32'h00000186;
      12'b001000101000 : romData <= 32'h04004186;
      12'b001000101001 : romData <= 32'h08008186;
      12'b001000101010 : romData <= 32'h0C00C186;
      12'b001000101011 : romData <= 32'h10000187;
      12'b001000101100 : romData <= 32'h14004187;
      12'b001000101101 : romData <= 32'h18002185;
      12'b001000101110 : romData <= 32'h00480044;
      12'b001000101111 : romData <= 32'h1C00219C;
      12'b001000110000 : romData <= 32'h0400169F;
      12'b001000110001 : romData <= 32'h04A074E0;
      12'b001000110010 : romData <= 32'h0000D686;
      12'b001000110011 : romData <= 32'h61FFFF07;
      12'b001000110100 : romData <= 32'h04B096E0;
      12'b001000110101 : romData <= 32'h0000201A;
      12'b001000110110 : romData <= 32'h008810E4;
      12'b001000110111 : romData <= 32'h04000010;
      12'b001000111000 : romData <= 32'h04B096E0;
      12'b001000111001 : romData <= 32'h5BFFFF07;
      12'b001000111010 : romData <= 32'h048070E0;
      12'b001000111011 : romData <= 32'h04C0D8E2;
      12'b001000111100 : romData <= 32'h0100529E;
      12'b001000111101 : romData <= 32'hABFFFF03;
      12'b001000111110 : romData <= 32'h0100529E;
      12'b001000111111 : romData <= 32'h00005686;
      12'b001001000000 : romData <= 32'h00A00048;
      12'b001001000001 : romData <= 32'h049072E0;
      12'b001001000010 : romData <= 32'h0000201A;
      12'b001001000011 : romData <= 32'h008810E4;
      12'b001001000100 : romData <= 32'hE3FFFF13;
      12'b001001000101 : romData <= 32'h049072E0;
      12'b001001000110 : romData <= 32'hDFFFFF03;
      12'b001001000111 : romData <= 32'h00000015;
      12'b001001001000 : romData <= 32'h00A00048;
      12'b001001001001 : romData <= 32'h04C078E0;
      12'b001001001010 : romData <= 32'h0000201A;
      12'b001001001011 : romData <= 32'h008810E4;
      12'b001001001100 : romData <= 32'hF1FFFF13;
      12'b001001001101 : romData <= 32'h00000015;
      12'b001001001110 : romData <= 32'h00800048;
      12'b001001001111 : romData <= 32'h04C078E0;
      12'b001001010000 : romData <= 32'h98FFFF03;
      12'b001001010001 : romData <= 32'h0100529E;
      12'b001001010010 : romData <= 32'h0050201A;
      12'b001001010011 : romData <= 32'h030071AA;
      12'b001001010100 : romData <= 32'h83FFA0AE;
      12'b001001010101 : romData <= 32'h00A813D8;
      12'b001001010110 : romData <= 32'h1B00A0AA;
      12'b001001010111 : romData <= 32'h00A811D8;
      12'b001001011000 : romData <= 32'h010031AA;
      12'b001001011001 : romData <= 32'h000011D8;
      12'b001001011010 : romData <= 32'h030020AA;
      12'b001001011011 : romData <= 32'h008813D8;
      12'b001001011100 : romData <= 32'h00480044;
      12'b001001011101 : romData <= 32'h00000015;
      12'b001001011110 : romData <= 32'h0050601A;
      12'b001001011111 : romData <= 32'h0500B3AA;
      12'b001001100000 : romData <= 32'h0000358E;
      12'b001001100001 : romData <= 32'h400031A6;
      12'b001001100010 : romData <= 32'h0000E01A;
      12'b001001100011 : romData <= 32'h00B811E4;
      12'b001001100100 : romData <= 32'h05000010;
      12'b001001100101 : romData <= 32'h00000015;
      12'b001001100110 : romData <= 32'h001813D8;
      12'b001001100111 : romData <= 32'h00480044;
      12'b001001101000 : romData <= 32'h00000015;
      12'b001001101001 : romData <= 32'h00000015;
      12'b001001101010 : romData <= 32'hF6FFFF03;
      12'b001001101011 : romData <= 32'h00000015;
      12'b001001101100 : romData <= 32'h0050601A;
      12'b001001101101 : romData <= 32'h0500B3AA;
      12'b001001101110 : romData <= 32'h0000358E;
      12'b001001101111 : romData <= 32'h010031A6;
      12'b001001110000 : romData <= 32'h0000E01A;
      12'b001001110001 : romData <= 32'h00B811E4;
      12'b001001110010 : romData <= 32'hFCFFFF13;
      12'b001001110011 : romData <= 32'h00000015;
      12'b001001110100 : romData <= 32'h0000738D;
      12'b001001110101 : romData <= 32'h00480044;
      12'b001001110110 : romData <= 32'h00000015;
      12'b001001110111 : romData <= 32'hF8FF219C;
      12'b001001111000 : romData <= 32'hFF0063A4;
      12'b001001111001 : romData <= 32'h008001D4;
      12'b001001111010 : romData <= 32'hD0FF039E;
      12'b001001111011 : romData <= 32'hFF0030A6;
      12'b001001111100 : romData <= 32'h090060AA;
      12'b001001111101 : romData <= 32'h009851E4;
      12'b001001111110 : romData <= 32'h0800000C;
      12'b001001111111 : romData <= 32'h044801D4;
      12'b001010000000 : romData <= 32'hBFFF239E;
      12'b001010000001 : romData <= 32'hFF0031A6;
      12'b001010000010 : romData <= 32'h050060AA;
      12'b001010000011 : romData <= 32'h009851E4;
      12'b001010000100 : romData <= 32'h12000010;
      12'b001010000101 : romData <= 32'hC9FF039E;
      12'b001010000110 : romData <= 32'hE6FFFF07;
      12'b001010000111 : romData <= 32'h00000015;
      12'b001010001000 : romData <= 32'hFF006BA5;
      12'b001010001001 : romData <= 32'hD0FF6B9E;
      12'b001010001010 : romData <= 32'hFF00B3A6;
      12'b001010001011 : romData <= 32'h0900E0AA;
      12'b001010001100 : romData <= 32'hBFFF2B9E;
      12'b001010001101 : romData <= 32'h00B855E4;
      12'b001010001110 : romData <= 32'h10000010;
      12'b001010001111 : romData <= 32'hFF0031A6;
      12'b001010010000 : romData <= 32'h040020AA;
      12'b001010010001 : romData <= 32'h088810E2;
      12'b001010010010 : romData <= 32'hF4FFFF03;
      12'b001010010011 : romData <= 32'h008013E2;
      12'b001010010100 : romData <= 32'hF2FFFF03;
      12'b001010010101 : romData <= 32'h0000001A;
      12'b001010010110 : romData <= 32'h9FFF239E;
      12'b001010010111 : romData <= 32'hFF0031A6;
      12'b001010011000 : romData <= 32'h050060AA;
      12'b001010011001 : romData <= 32'h009851E4;
      12'b001010011010 : romData <= 32'hFAFFFF13;
      12'b001010011011 : romData <= 32'h00000015;
      12'b001010011100 : romData <= 32'hEAFFFF03;
      12'b001010011101 : romData <= 32'hA9FF039E;
      12'b001010011110 : romData <= 32'h050060AA;
      12'b001010011111 : romData <= 32'h009851E4;
      12'b001010100000 : romData <= 32'h06000010;
      12'b001010100001 : romData <= 32'h040020AA;
      12'b001010100010 : romData <= 32'h088810E2;
      12'b001010100011 : romData <= 32'hC9FF6B9D;
      12'b001010100100 : romData <= 32'hE2FFFF03;
      12'b001010100101 : romData <= 32'h00800BE2;
      12'b001010100110 : romData <= 32'h9FFF2B9E;
      12'b001010100111 : romData <= 32'hFF0031A6;
      12'b001010101000 : romData <= 32'h050060AA;
      12'b001010101001 : romData <= 32'h009851E4;
      12'b001010101010 : romData <= 32'h05000010;
      12'b001010101011 : romData <= 32'h040020AA;
      12'b001010101100 : romData <= 32'h088810E2;
      12'b001010101101 : romData <= 32'hF7FFFF03;
      12'b001010101110 : romData <= 32'hA9FF6B9D;
      12'b001010101111 : romData <= 32'h048070E1;
      12'b001010110000 : romData <= 32'h04002185;
      12'b001010110001 : romData <= 32'h00000186;
      12'b001010110010 : romData <= 32'h00480044;
      12'b001010110011 : romData <= 32'h0800219C;
      12'b001010110100 : romData <= 32'hFF0063A4;
      12'b001010110101 : romData <= 32'h020020AA;
      12'b001010110110 : romData <= 32'h00191170;
      12'b001010110111 : romData <= 32'h00480044;
      12'b001010111000 : romData <= 32'h00000015;
      12'b001010111001 : romData <= 32'h041863E1;
      12'b001010111010 : romData <= 32'h0000201A;
      12'b001010111011 : romData <= 32'h002831E4;
      12'b001010111100 : romData <= 32'h04000010;
      12'b001010111101 : romData <= 32'h008864E2;
      12'b001010111110 : romData <= 32'h00480044;
      12'b001010111111 : romData <= 32'h00000015;
      12'b001011000000 : romData <= 32'h0000B392;
      12'b001011000001 : romData <= 32'h00886BE2;
      12'b001011000010 : romData <= 32'h00A813D8;
      12'b001011000011 : romData <= 32'hF8FFFF03;
      12'b001011000100 : romData <= 32'h0100319E;
      12'b001011000101 : romData <= 32'h0000201A;
      12'b001011000110 : romData <= 32'hFFFFE01A;
      12'b001011000111 : romData <= 32'h020060AA;
      12'b001011001000 : romData <= 32'h0898B1E2;
      12'b001011001001 : romData <= 32'h100060AA;
      12'b001011001010 : romData <= 32'h089871E2;
      12'b001011001011 : romData <= 32'h05B873E2;
      12'b001011001100 : romData <= 32'h048873E2;
      12'b001011001101 : romData <= 32'h009815D4;
      12'b001011001110 : romData <= 32'h0100319E;
      12'b001011001111 : romData <= 32'h002060AA;
      12'b001011010000 : romData <= 32'h009831E4;
      12'b001011010001 : romData <= 32'hF6FFFF13;
      12'b001011010010 : romData <= 32'h0000A01A;
      12'b001011010011 : romData <= 32'h0000201A;
      12'b001011010100 : romData <= 32'hFFFFE01A;
      12'b001011010101 : romData <= 32'h020060AA;
      12'b001011010110 : romData <= 32'h089871E2;
      12'b001011010111 : romData <= 32'h00003387;
      12'b001011011000 : romData <= 32'h100060AA;
      12'b001011011001 : romData <= 32'h089871E2;
      12'b001011011010 : romData <= 32'h05B873E2;
      12'b001011011011 : romData <= 32'h048873E2;
      12'b001011011100 : romData <= 32'h009819E4;
      12'b001011011101 : romData <= 32'h03000010;
      12'b001011011110 : romData <= 32'h00000015;
      12'b001011011111 : romData <= 32'h0100B59E;
      12'b001011100000 : romData <= 32'h0100319E;
      12'b001011100001 : romData <= 32'h002060AA;
      12'b001011100010 : romData <= 32'h009831E4;
      12'b001011100011 : romData <= 32'hF2FFFF13;
      12'b001011100100 : romData <= 32'h00000015;
      12'b001011100101 : romData <= 32'h0000201A;
      12'b001011100110 : romData <= 32'h008815E4;
      12'b001011100111 : romData <= 32'h54000010;
      12'b001011101000 : romData <= 32'h010020AA;
      12'b001011101001 : romData <= 32'h018860C3;
      12'b001011101010 : romData <= 32'h0000A01A;
      12'b001011101011 : romData <= 32'h0000201A;
      12'b001011101100 : romData <= 32'hFFFFE01A;
      12'b001011101101 : romData <= 32'h020060AA;
      12'b001011101110 : romData <= 32'h089871E2;
      12'b001011101111 : romData <= 32'h00003387;
      12'b001011110000 : romData <= 32'h100060AA;
      12'b001011110001 : romData <= 32'h089871E2;
      12'b001011110010 : romData <= 32'h05B873E2;
      12'b001011110011 : romData <= 32'h048873E2;
      12'b001011110100 : romData <= 32'h009819E4;
      12'b001011110101 : romData <= 32'h03000010;
      12'b001011110110 : romData <= 32'h00000015;
      12'b001011110111 : romData <= 32'h0100B59E;
      12'b001011111000 : romData <= 32'h0100319E;
      12'b001011111001 : romData <= 32'h002060AA;
      12'b001011111010 : romData <= 32'h009831E4;
      12'b001011111011 : romData <= 32'hF2FFFF13;
      12'b001011111100 : romData <= 32'h00000015;
      12'b001011111101 : romData <= 32'h0000201A;
      12'b001011111110 : romData <= 32'h008815E4;
      12'b001011111111 : romData <= 32'h3C000010;
      12'b001100000000 : romData <= 32'h020020AA;
      12'b001100000001 : romData <= 32'h018860C3;
      12'b001100000010 : romData <= 32'h0000A01A;
      12'b001100000011 : romData <= 32'h0000201A;
      12'b001100000100 : romData <= 32'hFFFFE01A;
      12'b001100000101 : romData <= 32'h020060AA;
      12'b001100000110 : romData <= 32'h089871E2;
      12'b001100000111 : romData <= 32'h00003387;
      12'b001100001000 : romData <= 32'h100060AA;
      12'b001100001001 : romData <= 32'h089871E2;
      12'b001100001010 : romData <= 32'h05B873E2;
      12'b001100001011 : romData <= 32'h048873E2;
      12'b001100001100 : romData <= 32'h009819E4;
      12'b001100001101 : romData <= 32'h03000010;
      12'b001100001110 : romData <= 32'h00000015;
      12'b001100001111 : romData <= 32'h0100B59E;
      12'b001100010000 : romData <= 32'h0100319E;
      12'b001100010001 : romData <= 32'h002060AA;
      12'b001100010010 : romData <= 32'h009831E4;
      12'b001100010011 : romData <= 32'hF2FFFF13;
      12'b001100010100 : romData <= 32'h00000015;
      12'b001100010101 : romData <= 32'h0000201A;
      12'b001100010110 : romData <= 32'h008815E4;
      12'b001100010111 : romData <= 32'h24000010;
      12'b001100011000 : romData <= 32'h030020AA;
      12'b001100011001 : romData <= 32'h018860C3;
      12'b001100011010 : romData <= 32'h0000A01A;
      12'b001100011011 : romData <= 32'h0000201A;
      12'b001100011100 : romData <= 32'hFFFFE01A;
      12'b001100011101 : romData <= 32'h020060AA;
      12'b001100011110 : romData <= 32'h089871E2;
      12'b001100011111 : romData <= 32'h00003387;
      12'b001100100000 : romData <= 32'h100060AA;
      12'b001100100001 : romData <= 32'h089871E2;
      12'b001100100010 : romData <= 32'h05B873E2;
      12'b001100100011 : romData <= 32'h048873E2;
      12'b001100100100 : romData <= 32'h009819E4;
      12'b001100100101 : romData <= 32'h03000010;
      12'b001100100110 : romData <= 32'h00000015;
      12'b001100100111 : romData <= 32'h0100B59E;
      12'b001100101000 : romData <= 32'h0100319E;
      12'b001100101001 : romData <= 32'h002060AA;
      12'b001100101010 : romData <= 32'h009831E4;
      12'b001100101011 : romData <= 32'hF2FFFF13;
      12'b001100101100 : romData <= 32'h00000015;
      12'b001100101101 : romData <= 32'h0000201A;
      12'b001100101110 : romData <= 32'h008815E4;
      12'b001100101111 : romData <= 32'h0C000010;
      12'b001100110000 : romData <= 32'h00F0A018;
      12'b001100110001 : romData <= 32'h00F08018;
      12'b001100110010 : romData <= 32'h00F06018;
      12'b001100110011 : romData <= 32'hFCFF219C;
      12'b001100110100 : romData <= 32'h271EA59C;
      12'b001100110101 : romData <= 32'h7809849C;
      12'b001100110110 : romData <= 32'h004801D4;
      12'b001100110111 : romData <= 32'hA4FEFF07;
      12'b001100111000 : romData <= 32'hD00A639C;
      12'b001100111010 : romData <= 32'h00000015;
      12'b001100111011 : romData <= 32'h00480044;
      12'b001100111100 : romData <= 32'h00000015;
      12'b001100111101 : romData <= 32'h9CFF219C;
      12'b001100111110 : romData <= 32'h00F08018;
      12'b001100111111 : romData <= 32'h3C00A0A8;
      12'b001101000000 : romData <= 32'hAC25849C;
      12'b001101000001 : romData <= 32'h508001D4;
      12'b001101000010 : romData <= 32'h549001D4;
      12'b001101000011 : romData <= 32'h58A001D4;
      12'b001101000100 : romData <= 32'h5CB001D4;
      12'b001101000101 : romData <= 32'h604801D4;
      12'b001101000110 : romData <= 32'h73FFFF07;
      12'b001101000111 : romData <= 32'h1400619C;
      12'b001101001000 : romData <= 32'h030020AA;
      12'b001101001001 : romData <= 32'h00011170;
      12'b001101001010 : romData <= 32'h090040B6;
      12'b001101001011 : romData <= 32'hFF0020AA;
      12'b001101001100 : romData <= 32'h0088B2E4;
      12'b001101001101 : romData <= 32'hFDFFFF13;
      12'b001101001110 : romData <= 32'h0F00D2A6;
      12'b001101001111 : romData <= 32'h010020AA;
      12'b001101010000 : romData <= 32'h008836E4;
      12'b001101010001 : romData <= 32'h34000010;
      12'b001101010010 : romData <= 32'h0000001A;
      12'b001101010011 : romData <= 32'h72FFFF07;
      12'b001101010100 : romData <= 32'h00000015;
      12'b001101010101 : romData <= 32'hADDE201A;
      12'b001101010110 : romData <= 32'h0004A01A;
      12'b001101010111 : romData <= 32'h001331AA;
      12'b001101011000 : romData <= 32'h00007586;
      12'b001101011001 : romData <= 32'h008833E4;
      12'b001101011010 : romData <= 32'h86000010;
      12'b001101011011 : romData <= 32'h00F0001A;
      12'b001101011100 : romData <= 32'h0050201A;
      12'b001101011101 : romData <= 32'h0200601A;
      12'b001101011110 : romData <= 32'h8C0031AA;
      12'b001101011111 : romData <= 32'h00003186;
      12'b001101100000 : romData <= 32'h039831E2;
      12'b001101100001 : romData <= 32'h0000601A;
      12'b001101100010 : romData <= 32'h009831E4;
      12'b001101100011 : romData <= 32'h22000010;
      12'b001101100100 : romData <= 32'h7809109E;
      12'b001101100101 : romData <= 32'h040075AA;
      12'b001101100110 : romData <= 32'h0200E0AA;
      12'b001101100111 : romData <= 32'h00007386;
      12'b001101101000 : romData <= 32'h08B873E2;
      12'b001101101001 : romData <= 32'h009831E4;
      12'b001101101010 : romData <= 32'h71000010;
      12'b001101101011 : romData <= 32'h0088F5E2;
      12'b001101101100 : romData <= 32'h00F0001A;
      12'b001101101101 : romData <= 32'h7809109E;
      12'b001101101110 : romData <= 32'h00F06018;
      12'b001101101111 : romData <= 32'h00F0A018;
      12'b001101110000 : romData <= 32'hD00A639C;
      12'b001101110001 : romData <= 32'h5B22A59C;
      12'b001101110010 : romData <= 32'h048090E0;
      12'b001101110011 : romData <= 32'h68FEFF07;
      12'b001101110100 : romData <= 32'h101801D4;
      12'b001101110101 : romData <= 32'h110080B6;
      12'b001101110110 : romData <= 32'hFFBF20AE;
      12'b001101110111 : romData <= 32'h038834E2;
      12'b001101111000 : romData <= 32'h118800C0;
      12'b001101111001 : romData <= 32'h0D0040AA;
      12'b001101111010 : romData <= 32'h00E052B6;
      12'b001101111011 : romData <= 32'h00F0A018;
      12'b001101111100 : romData <= 32'h009001D4;
      12'b001101111101 : romData <= 32'h5F1EA59C;
      12'b001101111110 : romData <= 32'h048090E0;
      12'b001101111111 : romData <= 32'h5CFEFF07;
      12'b001110000000 : romData <= 32'h10006184;
      12'b001110000001 : romData <= 32'hE7BF20AE;
      12'b001110000010 : romData <= 32'h038894E2;
      12'b001110000011 : romData <= 32'h00900044;
      12'b001110000100 : romData <= 32'h11A000C0;
      12'b001110000101 : romData <= 32'h00F0801A;
      12'b001110000110 : romData <= 32'hD00A949E;
      12'b001110000111 : romData <= 32'h00F0A018;
      12'b001110001000 : romData <= 32'h048090E0;
      12'b001110001001 : romData <= 32'h7A1EA59C;
      12'b001110001010 : romData <= 32'h51FEFF07;
      12'b001110001011 : romData <= 32'h04A074E0;
      12'b001110001100 : romData <= 32'h00F0A018;
      12'b001110001101 : romData <= 32'h048090E0;
      12'b001110001110 : romData <= 32'hA91EA59C;
      12'b001110001111 : romData <= 32'h4CFEFF07;
      12'b001110010000 : romData <= 32'h04A074E0;
      12'b001110010001 : romData <= 32'h00F0A018;
      12'b001110010010 : romData <= 32'h048090E0;
      12'b001110010011 : romData <= 32'hCC1EA59C;
      12'b001110010100 : romData <= 32'h47FEFF07;
      12'b001110010101 : romData <= 32'h04A074E0;
      12'b001110010110 : romData <= 32'h040020AA;
      12'b001110010111 : romData <= 32'h488832E2;
      12'b001110011000 : romData <= 32'h0F0031A6;
      12'b001110011001 : romData <= 32'h00F0A018;
      12'b001110011010 : romData <= 32'h048090E0;
      12'b001110011011 : romData <= 32'h048801D4;
      12'b001110011100 : romData <= 32'hFE1EA59C;
      12'b001110011101 : romData <= 32'h04A074E0;
      12'b001110011110 : romData <= 32'h3DFEFF07;
      12'b001110011111 : romData <= 32'h00B001D4;
      12'b001110100000 : romData <= 32'h0C0020AA;
      12'b001110100001 : romData <= 32'h488832E2;
      12'b001110100010 : romData <= 32'h0F0031A6;
      12'b001110100011 : romData <= 32'h0C8801D4;
      12'b001110100100 : romData <= 32'h100020AA;
      12'b001110100101 : romData <= 32'h488832E2;
      12'b001110100110 : romData <= 32'h0F0031A6;
      12'b001110100111 : romData <= 32'h088801D4;
      12'b001110101000 : romData <= 32'h140020AA;
      12'b001110101001 : romData <= 32'h488832E2;
      12'b001110101010 : romData <= 32'h0F0031A6;
      12'b001110101011 : romData <= 32'h048801D4;
      12'b001110101100 : romData <= 32'h180020AA;
      12'b001110101101 : romData <= 32'h488852E2;
      12'b001110101110 : romData <= 32'h0F0052A6;
      12'b001110101111 : romData <= 32'h00F0A018;
      12'b001110110000 : romData <= 32'h009001D4;
      12'b001110110001 : romData <= 32'h048090E0;
      12'b001110110010 : romData <= 32'h1C1FA59C;
      12'b001110110011 : romData <= 32'h04A074E0;
      12'b001110110100 : romData <= 32'h27FEFF07;
      12'b001110110101 : romData <= 32'h00F0401A;
      12'b001110110110 : romData <= 32'h1400019E;
      12'b001110110111 : romData <= 32'h7809529E;
      12'b001110111000 : romData <= 32'h0000201A;
      12'b001110111001 : romData <= 32'h0000B084;
      12'b001110111010 : romData <= 32'h008825E4;
      12'b001110111011 : romData <= 32'h27000010;
      12'b001110111100 : romData <= 32'h010020AA;
      12'b001110111101 : romData <= 32'h008836E4;
      12'b001110111110 : romData <= 32'h1600000C;
      12'b001110111111 : romData <= 32'h00000015;
      12'b001111000000 : romData <= 32'h00F0A018;
      12'b001111000001 : romData <= 32'h2D1FA59C;
      12'b001111000010 : romData <= 32'h00008018;
      12'b001111000011 : romData <= 32'h18FEFF07;
      12'b001111000100 : romData <= 32'h04A074E0;
      12'b001111000101 : romData <= 32'h025020B6;
      12'b001111000110 : romData <= 32'h0000601A;
      12'b001111000111 : romData <= 32'h009871E5;
      12'b001111001000 : romData <= 32'hFDFFFF13;
      12'b001111001001 : romData <= 32'h00000015;
      12'b001111001010 : romData <= 32'h035000B6;
      12'b001111001011 : romData <= 32'h00F0A018;
      12'b001111001100 : romData <= 32'h008001D4;
      12'b001111001101 : romData <= 32'h4F1FA59C;
      12'b001111001110 : romData <= 32'h00008018;
      12'b001111001111 : romData <= 32'h0CFEFF07;
      12'b001111010000 : romData <= 32'h04A074E0;
      12'b001111010001 : romData <= 32'h00800044;
      12'b001111010010 : romData <= 32'h00000015;
      12'b001111010011 : romData <= 32'h00000015;
      12'b001111010100 : romData <= 32'h50000186;
      12'b001111010101 : romData <= 32'h54004186;
      12'b001111010110 : romData <= 32'h58008186;
      12'b001111010111 : romData <= 32'h5C00C186;
      12'b001111011000 : romData <= 32'h60002185;
      12'b001111011001 : romData <= 32'h00480044;
      12'b001111011010 : romData <= 32'h6400219C;
      12'b001111011011 : romData <= 32'h0000F786;
      12'b001111011100 : romData <= 32'h0400319E;
      12'b001111011101 : romData <= 32'hFCBFF1D7;
      12'b001111011110 : romData <= 32'h8CFFFF03;
      12'b001111011111 : romData <= 32'h009831E4;
      12'b001111100000 : romData <= 32'hA5FFFF03;
      12'b001111100001 : romData <= 32'h7809109E;
      12'b001111100010 : romData <= 32'h008816E4;
      12'b001111100011 : romData <= 32'hDDFFFF0F;
      12'b001111100100 : romData <= 32'h049092E0;
      12'b001111100101 : romData <= 32'h04A074E0;
      12'b001111100110 : romData <= 32'hF5FDFF07;
      12'b001111100111 : romData <= 32'h0400109E;
      12'b001111101000 : romData <= 32'hD1FFFF03;
      12'b001111101001 : romData <= 32'h0000201A;
      12'b001111101010 : romData <= 32'hADDE201A;
      12'b001111101011 : romData <= 32'h001371AA;
      12'b001111101100 : romData <= 32'h009803E4;
      12'b001111101101 : romData <= 32'h14000010;
      12'b001111101110 : romData <= 32'h00006019;
      12'b001111101111 : romData <= 32'hFFFF601A;
      12'b001111110000 : romData <= 32'h039863E0;
      12'b001111110001 : romData <= 32'h008823E4;
      12'b001111110010 : romData <= 32'h0F000010;
      12'b001111110011 : romData <= 32'hFFFF60AD;
      12'b001111110100 : romData <= 32'h00F0A018;
      12'b001111110101 : romData <= 32'h00F08018;
      12'b001111110110 : romData <= 32'h00F06018;
      12'b001111110111 : romData <= 32'hFCFF219C;
      12'b001111111000 : romData <= 32'h6E1FA59C;
      12'b001111111001 : romData <= 32'h7809849C;
      12'b001111111010 : romData <= 32'h004801D4;
      12'b001111111011 : romData <= 32'hE0FDFF07;
      12'b001111111100 : romData <= 32'hD00A639C;
      12'b001111111101 : romData <= 32'hFFFF60AD;
      12'b001111111110 : romData <= 32'h00002185;
      12'b001111111111 : romData <= 32'h00480044;
      12'b010000000000 : romData <= 32'h0400219C;
      12'b010000000001 : romData <= 32'h00480044;
      12'b010000000010 : romData <= 32'h00000015;
      12'b010000000011 : romData <= 32'hACFC219C;
      12'b010000000100 : romData <= 32'h287301D4;
      12'b010000000101 : romData <= 32'h2C8301D4;
      12'b010000000110 : romData <= 32'h309301D4;
      12'b010000000111 : romData <= 32'h34A301D4;
      12'b010000001000 : romData <= 32'h38B301D4;
      12'b010000001001 : romData <= 32'h3CC301D4;
      12'b010000001010 : romData <= 32'h40D301D4;
      12'b010000001011 : romData <= 32'h44E301D4;
      12'b010000001100 : romData <= 32'h48F301D4;
      12'b010000001101 : romData <= 32'h4C1301D4;
      12'b010000001110 : romData <= 32'h504B01D4;
      12'b010000001111 : romData <= 32'h00C0201A;
      12'b010000010000 : romData <= 32'h068800C0;
      12'b010000010001 : romData <= 32'h110020B6;
      12'b010000010010 : romData <= 32'h248801D4;
      12'b010000010011 : romData <= 32'h24002186;
      12'b010000010100 : romData <= 32'h100031AA;
      12'b010000010101 : romData <= 32'h248801D4;
      12'b010000010110 : romData <= 32'h24002186;
      12'b010000010111 : romData <= 32'h118800C0;
      12'b010000011000 : romData <= 32'h3AFEFF07;
      12'b010000011001 : romData <= 32'h7F00C019;
      12'b010000011010 : romData <= 32'h23FFFF07;
      12'b010000011011 : romData <= 32'h010040AA;
      12'b010000011100 : romData <= 32'h00F0201A;
      12'b010000011101 : romData <= 32'h6C22319E;
      12'b010000011110 : romData <= 32'hFCFFCEA9;
      12'b010000011111 : romData <= 32'h0000C01B;
      12'b010000100000 : romData <= 32'h0000001B;
      12'b010000100001 : romData <= 32'h049052E0;
      12'b010000100010 : romData <= 32'h0000001A;
      12'b010000100011 : romData <= 32'h148801D4;
      12'b010000100100 : romData <= 32'h48FEFF07;
      12'b010000100101 : romData <= 32'h00000015;
      12'b010000100110 : romData <= 32'hFF002BA6;
      12'b010000100111 : romData <= 32'h270060AA;
      12'b010000101000 : romData <= 32'h009811E4;
      12'b010000101001 : romData <= 32'hA0020010;
      12'b010000101010 : romData <= 32'h04584BE3;
      12'b010000101011 : romData <= 32'h009851E4;
      12'b010000101100 : romData <= 32'h47000010;
      12'b010000101101 : romData <= 32'h230060AA;
      12'b010000101110 : romData <= 32'h009811E4;
      12'b010000101111 : romData <= 32'h87000010;
      12'b010000110000 : romData <= 32'h009851E4;
      12'b010000110001 : romData <= 32'h10000010;
      12'b010000110010 : romData <= 32'h160060AA;
      12'b010000110011 : romData <= 32'hF6FF319E;
      12'b010000110100 : romData <= 32'hFF0031A6;
      12'b010000110101 : romData <= 32'h009851E4;
      12'b010000110110 : romData <= 32'h09000010;
      12'b010000110111 : romData <= 32'h4000601A;
      12'b010000111000 : romData <= 32'h090073AA;
      12'b010000111001 : romData <= 32'h488833E2;
      12'b010000111010 : romData <= 32'h010031A6;
      12'b010000111011 : romData <= 32'h0000601A;
      12'b010000111100 : romData <= 32'h009831E4;
      12'b010000111101 : romData <= 32'hE7FFFF13;
      12'b010000111110 : romData <= 32'h00000015;
      12'b010000111111 : romData <= 32'h45000000;
      12'b010001000000 : romData <= 32'h00006019;
      12'b010001000001 : romData <= 32'h260060AA;
      12'b010001000010 : romData <= 32'h009811E4;
      12'b010001000011 : romData <= 32'h4100000C;
      12'b010001000100 : romData <= 32'h00006019;
      12'b010001000101 : romData <= 32'h27FEFF07;
      12'b010001000110 : romData <= 32'h00000015;
      12'b010001000111 : romData <= 32'h00F0A018;
      12'b010001001000 : romData <= 32'h00F06018;
      12'b010001001001 : romData <= 32'hD01FA59C;
      12'b010001001010 : romData <= 32'h00008018;
      12'b010001001011 : romData <= 32'hD00A639C;
      12'b010001001100 : romData <= 32'h8FFDFF07;
      12'b010001001101 : romData <= 32'hFF004BA7;
      12'b010001001110 : romData <= 32'h0000201A;
      12'b010001001111 : romData <= 32'h200060AA;
      12'b010001010000 : romData <= 32'h00981AE4;
      12'b010001010001 : romData <= 32'h1D000010;
      12'b010001010010 : romData <= 32'h2800619E;
      12'b010001010011 : romData <= 32'h008891E3;
      12'b010001010100 : romData <= 32'h00889CE3;
      12'b010001010101 : romData <= 32'h0098BCE2;
      12'b010001010110 : romData <= 32'h0000601A;
      12'b010001010111 : romData <= 32'h0100739E;
      12'b010001011000 : romData <= 32'h00D015D8;
      12'b010001011001 : romData <= 32'h188801D4;
      12'b010001011010 : romData <= 32'h109801D4;
      12'b010001011011 : romData <= 32'h11FEFF07;
      12'b010001011100 : romData <= 32'h0CA801D4;
      12'b010001011101 : romData <= 32'h200020AA;
      12'b010001011110 : romData <= 32'hFF004BA7;
      12'b010001011111 : romData <= 32'h00883AE4;
      12'b010001100000 : romData <= 32'h0C00A186;
      12'b010001100001 : romData <= 32'h10006186;
      12'b010001100010 : romData <= 32'h0100B59E;
      12'b010001100011 : romData <= 32'hF4FFFF13;
      12'b010001100100 : romData <= 32'h18002186;
      12'b010001100101 : romData <= 32'h1003BC9E;
      12'b010001100110 : romData <= 32'h1800E19E;
      12'b010001100111 : romData <= 32'h00B895E3;
      12'b010001101000 : romData <= 32'h00989CE3;
      12'b010001101001 : romData <= 32'h0100319E;
      12'b010001101010 : romData <= 32'hFF0060AA;
      12'b010001101011 : romData <= 32'h0098B1E5;
      12'b010001101100 : romData <= 32'hB8FFFF0F;
      12'b010001101101 : romData <= 32'h0005FCDB;
      12'b010001101110 : romData <= 32'hFEFDFF07;
      12'b010001101111 : romData <= 32'h0C8801D4;
      12'b010001110000 : romData <= 32'hFF004BA7;
      12'b010001110001 : romData <= 32'hDEFFFF03;
      12'b010001110010 : romData <= 32'h0C002186;
      12'b010001110011 : romData <= 32'h2D0060AA;
      12'b010001110100 : romData <= 32'h009811E4;
      12'b010001110101 : romData <= 32'h0A000010;
      12'b010001110110 : romData <= 32'h009851E4;
      12'b010001110111 : romData <= 32'h24000010;
      12'b010001111000 : romData <= 32'h2A0060AA;
      12'b010001111001 : romData <= 32'h009811E4;
      12'b010001111010 : romData <= 32'h43000010;
      12'b010001111011 : romData <= 32'h2B0060AA;
      12'b010001111100 : romData <= 32'h009811E4;
      12'b010001111101 : romData <= 32'h0700000C;
      12'b010001111110 : romData <= 32'h00006019;
      12'b010001111111 : romData <= 32'hEDFDFF07;
      12'b010010000000 : romData <= 32'h00000015;
      12'b010010000001 : romData <= 32'h180020AA;
      12'b010010000010 : romData <= 32'h08886BE1;
      12'b010010000011 : romData <= 32'h88886BE1;
      12'b010010000100 : romData <= 32'h180060AA;
      12'b010010000101 : romData <= 32'h08983AE2;
      12'b010010000110 : romData <= 32'h889831E2;
      12'b010010000111 : romData <= 32'h2800A19E;
      12'b010010001000 : romData <= 32'h0000801B;
      12'b010010001001 : romData <= 32'h0000F592;
      12'b010010001010 : romData <= 32'h008837E4;
      12'b010010001011 : romData <= 32'h4B020010;
      12'b010010001100 : romData <= 32'h00000015;
      12'b010010001101 : romData <= 32'h0100F592;
      12'b010010001110 : romData <= 32'h005817E4;
      12'b010010001111 : romData <= 32'h4702000C;
      12'b010010010000 : romData <= 32'h00F0401B;
      12'b010010010001 : romData <= 32'h00F0201A;
      12'b010010010010 : romData <= 32'h4D23319E;
      12'b010010010011 : romData <= 32'h00405AAB;
      12'b010010010100 : romData <= 32'h0C8801D4;
      12'b010010010101 : romData <= 32'h0000201A;
      12'b010010010110 : romData <= 32'h008832E4;
      12'b010010010111 : romData <= 32'h48020010;
      12'b010010011000 : romData <= 32'h00000015;
      12'b010010011001 : romData <= 32'h8BFFFF03;
      12'b010010011010 : romData <= 32'h010040AA;
      12'b010010011011 : romData <= 32'h3D0060AA;
      12'b010010011100 : romData <= 32'h009811E4;
      12'b010010011101 : romData <= 32'hE2FFFF13;
      12'b010010011110 : romData <= 32'h400060AA;
      12'b010010011111 : romData <= 32'h009811E4;
      12'b010010100000 : romData <= 32'hE4FFFF0F;
      12'b010010100001 : romData <= 32'h00006019;
      12'b010010100010 : romData <= 32'hD5FDFF07;
      12'b010010100011 : romData <= 32'h200060A8;
      12'b010010100100 : romData <= 32'h080020AA;
      12'b010010100101 : romData <= 32'h00F0A018;
      12'b010010100110 : romData <= 32'h00F06018;
      12'b010010100111 : romData <= 32'h08888BE2;
      12'b010010101000 : romData <= 32'h005801D4;
      12'b010010101001 : romData <= 32'h0A0020AA;
      12'b010010101010 : romData <= 32'hE41FA59C;
      12'b010010101011 : romData <= 32'h00008018;
      12'b010010101100 : romData <= 32'hD00A639C;
      12'b010010101101 : romData <= 32'h488894E2;
      12'b010010101110 : romData <= 32'h2DFDFF07;
      12'b010010101111 : romData <= 32'h0458CBE2;
      12'b010010110000 : romData <= 32'h0000201A;
      12'b010010110001 : romData <= 32'h008814E4;
      12'b010010110010 : romData <= 32'h88020010;
      12'b010010110011 : romData <= 32'h0000C01B;
      12'b010010110100 : romData <= 32'h70FFFF03;
      12'b010010110101 : romData <= 32'h00000015;
      12'b010010110110 : romData <= 32'h00F0A018;
      12'b010010110111 : romData <= 32'hC01FA59C;
      12'b010010111000 : romData <= 32'h00F08018;
      12'b010010111001 : romData <= 32'h7809849C;
      12'b010010111010 : romData <= 32'h00F06018;
      12'b010010111011 : romData <= 32'h2D010000;
      12'b010010111100 : romData <= 32'hD00A639C;
      12'b010010111101 : romData <= 32'hAFFDFF07;
      12'b010010111110 : romData <= 32'h00000015;
      12'b010010111111 : romData <= 32'hFF006BA5;
      12'b010011000000 : romData <= 32'h6D0020AA;
      12'b010011000001 : romData <= 32'h00880BE4;
      12'b010011000010 : romData <= 32'h96010010;
      12'b010011000011 : romData <= 32'h00884BE4;
      12'b010011000100 : romData <= 32'h33000010;
      12'b010011000101 : romData <= 32'h660020AA;
      12'b010011000110 : romData <= 32'h00880BE4;
      12'b010011000111 : romData <= 32'h11010010;
      12'b010011001000 : romData <= 32'h00884BE4;
      12'b010011001001 : romData <= 32'h14000010;
      12'b010011001010 : romData <= 32'h630020AA;
      12'b010011001011 : romData <= 32'h00880BE4;
      12'b010011001100 : romData <= 32'hC9000010;
      12'b010011001101 : romData <= 32'h650020AA;
      12'b010011001110 : romData <= 32'h00880BE4;
      12'b010011001111 : romData <= 32'h60010010;
      12'b010011010000 : romData <= 32'h2A0020AA;
      12'b010011010001 : romData <= 32'h00880BE4;
      12'b010011010010 : romData <= 32'h52FFFF0F;
      12'b010011010011 : romData <= 32'h00000015;
      12'b010011010100 : romData <= 32'h00007084;
      12'b010011010101 : romData <= 32'h15FFFF07;
      12'b010011010110 : romData <= 32'h00000015;
      12'b010011010111 : romData <= 32'h0000201A;
      12'b010011011000 : romData <= 32'h00880BE4;
      12'b010011011001 : romData <= 32'h44000010;
      12'b010011011010 : romData <= 32'h00F0A018;
      12'b010011011011 : romData <= 32'hDDFFFF03;
      12'b010011011100 : romData <= 32'h0220A59C;
      12'b010011011101 : romData <= 32'h680020AA;
      12'b010011011110 : romData <= 32'h00880BE4;
      12'b010011011111 : romData <= 32'h62000010;
      12'b010011100000 : romData <= 32'h690020AA;
      12'b010011100001 : romData <= 32'h00880BE4;
      12'b010011100010 : romData <= 32'h42FFFF0F;
      12'b010011100011 : romData <= 32'h00000015;
      12'b010011100100 : romData <= 32'h00007084;
      12'b010011100101 : romData <= 32'h05FFFF07;
      12'b010011100110 : romData <= 32'h00000015;
      12'b010011100111 : romData <= 32'h0000201A;
      12'b010011101000 : romData <= 32'h00880BE4;
      12'b010011101001 : romData <= 32'h00F08018;
      12'b010011101010 : romData <= 32'h00F06018;
      12'b010011101011 : romData <= 32'h04003086;
      12'b010011101100 : romData <= 32'h7809849C;
      12'b010011101101 : romData <= 32'h81000010;
      12'b010011101110 : romData <= 32'hD00A639C;
      12'b010011101111 : romData <= 32'h00F0A018;
      12'b010011110000 : romData <= 32'h048801D4;
      12'b010011110001 : romData <= 32'h000001D4;
      12'b010011110010 : romData <= 32'h7820A59C;
      12'b010011110011 : romData <= 32'hE8FCFF07;
      12'b010011110100 : romData <= 32'h00000015;
      12'b010011110101 : romData <= 32'h2FFFFF03;
      12'b010011110110 : romData <= 32'h00000015;
      12'b010011110111 : romData <= 32'h730020AA;
      12'b010011111000 : romData <= 32'h00880BE4;
      12'b010011111001 : romData <= 32'h52000010;
      12'b010011111010 : romData <= 32'h00884BE4;
      12'b010011111011 : romData <= 32'h13000010;
      12'b010011111100 : romData <= 32'h710020AA;
      12'b010011111101 : romData <= 32'h00880BE4;
      12'b010011111110 : romData <= 32'hB8010010;
      12'b010011111111 : romData <= 32'h720020AA;
      12'b010100000000 : romData <= 32'h00880BE4;
      12'b010100000001 : romData <= 32'h4E000010;
      12'b010100000010 : romData <= 32'h700020AA;
      12'b010100000011 : romData <= 32'h00880BE4;
      12'b010100000100 : romData <= 32'h20FFFF0F;
      12'b010100000101 : romData <= 32'h00F0A018;
      12'b010100000110 : romData <= 32'h00F08018;
      12'b010100000111 : romData <= 32'h00F06018;
      12'b010100001000 : romData <= 32'h4F20A59C;
      12'b010100001001 : romData <= 32'h7809849C;
      12'b010100001010 : romData <= 32'hD1FCFF07;
      12'b010100001011 : romData <= 32'hD00A639C;
      12'b010100001100 : romData <= 32'h18FFFF03;
      12'b010100001101 : romData <= 32'h010040A8;
      12'b010100001110 : romData <= 32'h740020AA;
      12'b010100001111 : romData <= 32'h00880BE4;
      12'b010100010000 : romData <= 32'h67000010;
      12'b010100010001 : romData <= 32'h760020AA;
      12'b010100010010 : romData <= 32'h00880BE4;
      12'b010100010011 : romData <= 32'h11FFFF0F;
      12'b010100010100 : romData <= 32'h00F0A018;
      12'b010100010101 : romData <= 32'h00F08018;
      12'b010100010110 : romData <= 32'h00F06018;
      12'b010100010111 : romData <= 32'h6320A59C;
      12'b010100011000 : romData <= 32'h7809849C;
      12'b010100011001 : romData <= 32'hC2FCFF07;
      12'b010100011010 : romData <= 32'hD00A639C;
      12'b010100011011 : romData <= 32'h09FFFF03;
      12'b010100011100 : romData <= 32'h00004018;
      12'b010100011101 : romData <= 32'h00F0201A;
      12'b010100011110 : romData <= 32'h004031AA;
      12'b010100011111 : romData <= 32'h008830E4;
      12'b010100100000 : romData <= 32'h05000010;
      12'b010100100001 : romData <= 32'h010020AA;
      12'b010100100010 : romData <= 32'h0F8880C3;
      12'b010100100011 : romData <= 32'h01FFFF03;
      12'b010100100100 : romData <= 32'h00000015;
      12'b010100100101 : romData <= 32'h110020B6;
      12'b010100100110 : romData <= 32'hFFBF60AE;
      12'b010100100111 : romData <= 32'h248801D4;
      12'b010100101000 : romData <= 32'h24002186;
      12'b010100101001 : romData <= 32'h039831E2;
      12'b010100101010 : romData <= 32'h248801D4;
      12'b010100101011 : romData <= 32'h207040C1;
      12'b010100101100 : romData <= 32'h24002186;
      12'b010100101101 : romData <= 32'h118800C0;
      12'b010100101110 : romData <= 32'hE7BF60AE;
      12'b010100101111 : romData <= 32'h24002186;
      12'b010100110000 : romData <= 32'h039831E2;
      12'b010100110001 : romData <= 32'h248801D4;
      12'b010100110010 : romData <= 32'h0D0040AB;
      12'b010100110011 : romData <= 32'h00E05AB7;
      12'b010100110100 : romData <= 32'h00F0A018;
      12'b010100110101 : romData <= 32'h00F08018;
      12'b010100110110 : romData <= 32'h00F06018;
      12'b010100110111 : romData <= 32'h1D20A59C;
      12'b010100111000 : romData <= 32'h7809849C;
      12'b010100111001 : romData <= 32'hA2FCFF07;
      12'b010100111010 : romData <= 32'hD00A639C;
      12'b010100111011 : romData <= 32'h04D050E3;
      12'b010100111100 : romData <= 32'h24002186;
      12'b010100111101 : romData <= 32'h00D00044;
      12'b010100111110 : romData <= 32'h118800C0;
      12'b010100111111 : romData <= 32'hE5FEFF03;
      12'b010101000000 : romData <= 32'h00000015;
      12'b010101000001 : romData <= 32'h00F0A018;
      12'b010101000010 : romData <= 32'h00F06018;
      12'b010101000011 : romData <= 32'h2D22A59C;
      12'b010101000100 : romData <= 32'h00008018;
      12'b010101000101 : romData <= 32'h96FCFF07;
      12'b010101000110 : romData <= 32'h7809639C;
      12'b010101000111 : romData <= 32'hF6FDFF07;
      12'b010101001000 : romData <= 32'h00000015;
      12'b010101001001 : romData <= 32'hDBFEFF03;
      12'b010101001010 : romData <= 32'h00000015;
      12'b010101001011 : romData <= 32'hC8FBFF07;
      12'b010101001100 : romData <= 32'h00000015;
      12'b010101001101 : romData <= 32'hD7FEFF03;
      12'b010101001110 : romData <= 32'h00000015;
      12'b010101001111 : romData <= 32'h0004401B;
      12'b010101010000 : romData <= 32'h00007A84;
      12'b010101010001 : romData <= 32'h99FEFF07;
      12'b010101010010 : romData <= 32'h00000015;
      12'b010101010011 : romData <= 32'h0000201A;
      12'b010101010100 : romData <= 32'h00880BE4;
      12'b010101010101 : romData <= 32'h04000010;
      12'b010101010110 : romData <= 32'h00F0A018;
      12'b010101010111 : romData <= 32'h61FFFF03;
      12'b010101011000 : romData <= 32'h3220A59C;
      12'b010101011001 : romData <= 32'h04003AAA;
      12'b010101011010 : romData <= 32'h00007186;
      12'b010101011011 : romData <= 32'h020020AA;
      12'b010101011100 : romData <= 32'h088873E2;
      12'b010101011101 : romData <= 32'h0000201A;
      12'b010101011110 : romData <= 32'h009831E4;
      12'b010101011111 : romData <= 32'h0A000010;
      12'b010101100000 : romData <= 32'h0088BAE2;
      12'b010101100001 : romData <= 32'h110020B6;
      12'b010101100010 : romData <= 32'hFFBF60AE;
      12'b010101100011 : romData <= 32'h248801D4;
      12'b010101100100 : romData <= 32'h24002186;
      12'b010101100101 : romData <= 32'h039831E2;
      12'b010101100110 : romData <= 32'h248801D4;
      12'b010101100111 : romData <= 32'hC5FFFF03;
      12'b010101101000 : romData <= 32'h00000015;
      12'b010101101001 : romData <= 32'h0000B586;
      12'b010101101010 : romData <= 32'h0400319E;
      12'b010101101011 : romData <= 32'hFCAFF1D7;
      12'b010101101100 : romData <= 32'hF3FFFF03;
      12'b010101101101 : romData <= 32'h009831E4;
      12'b010101101110 : romData <= 32'h020060AA;
      12'b010101101111 : romData <= 32'h089831E2;
      12'b010101110000 : romData <= 32'h048031E2;
      12'b010101110001 : romData <= 32'hFFFF319E;
      12'b010101110010 : romData <= 32'h00F0A018;
      12'b010101110011 : romData <= 32'h048801D4;
      12'b010101110100 : romData <= 32'h008001D4;
      12'b010101110101 : romData <= 32'h7EFFFF03;
      12'b010101110110 : romData <= 32'h8C20A59C;
      12'b010101110111 : romData <= 32'h0000201A;
      12'b010101111000 : romData <= 32'h00F08018;
      12'b010101111001 : romData <= 32'h00F06018;
      12'b010101111010 : romData <= 32'h008830E4;
      12'b010101111011 : romData <= 32'h7809849C;
      12'b010101111100 : romData <= 32'h09000010;
      12'b010101111101 : romData <= 32'hD00A639C;
      12'b010101111110 : romData <= 32'h00F0A018;
      12'b010101111111 : romData <= 32'hAE20A59C;
      12'b010110000000 : romData <= 32'h5BFCFF07;
      12'b010110000001 : romData <= 32'h00F0001A;
      12'b010110000010 : romData <= 32'h0000001B;
      12'b010110000011 : romData <= 32'hA1FEFF03;
      12'b010110000100 : romData <= 32'h004010AA;
      12'b010110000101 : romData <= 32'h00F0201A;
      12'b010110000110 : romData <= 32'h004031AA;
      12'b010110000111 : romData <= 32'h008830E4;
      12'b010110001000 : romData <= 32'h08000010;
      12'b010110001001 : romData <= 32'h00F0A018;
      12'b010110001010 : romData <= 32'h00F0A018;
      12'b010110001011 : romData <= 32'h50FCFF07;
      12'b010110001100 : romData <= 32'hC520A59C;
      12'b010110001101 : romData <= 32'h0000001B;
      12'b010110001110 : romData <= 32'h96FEFF03;
      12'b010110001111 : romData <= 32'h0004001A;
      12'b010110010000 : romData <= 32'h4BFCFF07;
      12'b010110010001 : romData <= 32'hD820A59C;
      12'b010110010010 : romData <= 32'h0000001B;
      12'b010110010011 : romData <= 32'h91FEFF03;
      12'b010110010100 : romData <= 32'h0000001A;
      12'b010110010101 : romData <= 32'h00F0201A;
      12'b010110010110 : romData <= 32'h004031AA;
      12'b010110010111 : romData <= 32'h008810E4;
      12'b010110011000 : romData <= 32'h05000010;
      12'b010110011001 : romData <= 32'h0004201A;
      12'b010110011010 : romData <= 32'h008830E4;
      12'b010110011011 : romData <= 32'h05000010;
      12'b010110011100 : romData <= 32'h00000015;
      12'b010110011101 : romData <= 32'h00F0A018;
      12'b010110011110 : romData <= 32'h1AFFFF03;
      12'b010110011111 : romData <= 32'hEB20A59C;
      12'b010110100000 : romData <= 32'h00007084;
      12'b010110100001 : romData <= 32'h49FEFF07;
      12'b010110100010 : romData <= 32'h00000015;
      12'b010110100011 : romData <= 32'h0000201A;
      12'b010110100100 : romData <= 32'h00880BE4;
      12'b010110100101 : romData <= 32'h04000010;
      12'b010110100110 : romData <= 32'h00F0A018;
      12'b010110100111 : romData <= 32'h11FFFF03;
      12'b010110101000 : romData <= 32'h0D21A59C;
      12'b010110101001 : romData <= 32'h3F00201A;
      12'b010110101010 : romData <= 32'hFFFF31AA;
      12'b010110101011 : romData <= 32'h04007086;
      12'b010110101100 : romData <= 32'h0088B3E4;
      12'b010110101101 : romData <= 32'h23000010;
      12'b010110101110 : romData <= 32'h00F0A018;
      12'b010110101111 : romData <= 32'h09FFFF03;
      12'b010110110000 : romData <= 32'h2A21A59C;
      12'b010110110001 : romData <= 32'h0004201A;
      12'b010110110010 : romData <= 32'h0088BAE2;
      12'b010110110011 : romData <= 32'h00007587;
      12'b010110110100 : romData <= 32'h00003A87;
      12'b010110110101 : romData <= 32'h00C81BE4;
      12'b010110110110 : romData <= 32'h11000010;
      12'b010110110111 : romData <= 32'h04883AE2;
      12'b010110111000 : romData <= 32'h00F06018;
      12'b010110111001 : romData <= 32'h0000B586;
      12'b010110111010 : romData <= 32'h04E09CE0;
      12'b010110111011 : romData <= 32'h00003A87;
      12'b010110111100 : romData <= 32'hD00A639C;
      12'b010110111101 : romData <= 32'h08C801D4;
      12'b010110111110 : romData <= 32'h04A801D4;
      12'b010110111111 : romData <= 32'h008801D4;
      12'b010111000000 : romData <= 32'h18B801D4;
      12'b010111000001 : romData <= 32'h109801D4;
      12'b010111000010 : romData <= 32'h19FCFF07;
      12'b010111000011 : romData <= 32'h0C2801D4;
      12'b010111000100 : romData <= 32'h1800E186;
      12'b010111000101 : romData <= 32'h10006186;
      12'b010111000110 : romData <= 32'h0C00A184;
      12'b010111000111 : romData <= 32'h0100739E;
      12'b010111001000 : romData <= 32'h04005A9F;
      12'b010111001001 : romData <= 32'h00003786;
      12'b010111001010 : romData <= 32'h009851E4;
      12'b010111001011 : romData <= 32'hE6FFFF13;
      12'b010111001100 : romData <= 32'h00000015;
      12'b010111001101 : romData <= 32'h00F0A018;
      12'b010111001110 : romData <= 32'hEAFEFF03;
      12'b010111001111 : romData <= 32'h7021A59C;
      12'b010111010000 : romData <= 32'h00F0A018;
      12'b010111010001 : romData <= 32'h00F0801B;
      12'b010111010010 : romData <= 32'h0000401B;
      12'b010111010011 : romData <= 32'h0000601A;
      12'b010111010100 : romData <= 32'h0400E0AA;
      12'b010111010101 : romData <= 32'h4A21A59C;
      12'b010111010110 : romData <= 32'hF3FFFF03;
      12'b010111010111 : romData <= 32'h78099C9F;
      12'b010111011000 : romData <= 32'h00F0201A;
      12'b010111011001 : romData <= 32'h004031AA;
      12'b010111011010 : romData <= 32'h00F0801B;
      12'b010111011011 : romData <= 32'h00F0401B;
      12'b010111011100 : romData <= 32'h008810E4;
      12'b010111011101 : romData <= 32'h78099C9F;
      12'b010111011110 : romData <= 32'h06000010;
      12'b010111011111 : romData <= 32'hD00A5A9F;
      12'b010111100000 : romData <= 32'h0004201A;
      12'b010111100001 : romData <= 32'h008830E4;
      12'b010111100010 : romData <= 32'h0A000010;
      12'b010111100011 : romData <= 32'h00000015;
      12'b010111100100 : romData <= 32'h00F0A018;
      12'b010111100101 : romData <= 32'hEB20A59C;
      12'b010111100110 : romData <= 32'h04E09CE0;
      12'b010111100111 : romData <= 32'h04D07AE0;
      12'b010111101000 : romData <= 32'hF3FBFF07;
      12'b010111101001 : romData <= 32'h00000015;
      12'b010111101010 : romData <= 32'h3AFEFF03;
      12'b010111101011 : romData <= 32'h00000015;
      12'b010111101100 : romData <= 32'h00007084;
      12'b010111101101 : romData <= 32'hFDFDFF07;
      12'b010111101110 : romData <= 32'h00000015;
      12'b010111101111 : romData <= 32'h0000201A;
      12'b010111110000 : romData <= 32'h00880BE4;
      12'b010111110001 : romData <= 32'h04000010;
      12'b010111110010 : romData <= 32'h00F0A018;
      12'b010111110011 : romData <= 32'hF3FFFF03;
      12'b010111110100 : romData <= 32'h0D21A59C;
      12'b010111110101 : romData <= 32'h3F00201A;
      12'b010111110110 : romData <= 32'hFFFF31AA;
      12'b010111110111 : romData <= 32'h04007086;
      12'b010111111000 : romData <= 32'h0088B3E4;
      12'b010111111001 : romData <= 32'h04000010;
      12'b010111111010 : romData <= 32'h00F0A018;
      12'b010111111011 : romData <= 32'hEBFFFF03;
      12'b010111111100 : romData <= 32'h2A21A59C;
      12'b010111111101 : romData <= 32'h00F0A018;
      12'b010111111110 : romData <= 32'h7E21A59C;
      12'b010111111111 : romData <= 32'h04E09CE0;
      12'b011000000000 : romData <= 32'hDBFBFF07;
      12'b011000000001 : romData <= 32'h04D07AE0;
      12'b011000000010 : romData <= 32'h00F0A018;
      12'b011000000011 : romData <= 32'h0004201A;
      12'b011000000100 : romData <= 32'h0000601A;
      12'b011000000101 : romData <= 32'h00FCE01A;
      12'b011000000110 : romData <= 32'hA121A59C;
      12'b011000000111 : romData <= 32'h0400A0AA;
      12'b011000001000 : romData <= 32'h0000B586;
      12'b011000001001 : romData <= 32'h009855E4;
      12'b011000001010 : romData <= 32'h0F000010;
      12'b011000001011 : romData <= 32'hFFFF20AF;
      12'b011000001100 : romData <= 32'h00F0A018;
      12'b011000001101 : romData <= 32'hC821A59C;
      12'b011000001110 : romData <= 32'h04E09CE0;
      12'b011000001111 : romData <= 32'hCCFBFF07;
      12'b011000010000 : romData <= 32'h04D07AE0;
      12'b011000010001 : romData <= 32'h040020AA;
      12'b011000010010 : romData <= 32'h00006018;
      12'b011000010011 : romData <= 32'h00009184;
      12'b011000010100 : romData <= 32'hD5FAFF07;
      12'b011000010101 : romData <= 32'h00000015;
      12'b011000010110 : romData <= 32'h00F0A018;
      12'b011000010111 : romData <= 32'hCFFFFF03;
      12'b011000011000 : romData <= 32'hE121A59C;
      12'b011000011001 : romData <= 32'h0000B186;
      12'b011000011010 : romData <= 32'h00C815E4;
      12'b011000011011 : romData <= 32'h11000010;
      12'b011000011100 : romData <= 32'h00B8B1E2;
      12'b011000011101 : romData <= 32'h00A801D4;
      12'b011000011110 : romData <= 32'h04E09CE0;
      12'b011000011111 : romData <= 32'h04D07AE0;
      12'b011000100000 : romData <= 32'h209801D4;
      12'b011000100001 : romData <= 32'h1CB801D4;
      12'b011000100010 : romData <= 32'h188801D4;
      12'b011000100011 : romData <= 32'h0C2801D4;
      12'b011000100100 : romData <= 32'hB7FBFF07;
      12'b011000100101 : romData <= 32'h10A801D4;
      12'b011000100110 : romData <= 32'hBCFAFF07;
      12'b011000100111 : romData <= 32'h10006184;
      12'b011000101000 : romData <= 32'h20006186;
      12'b011000101001 : romData <= 32'h1C00E186;
      12'b011000101010 : romData <= 32'h18002186;
      12'b011000101011 : romData <= 32'h0C00A184;
      12'b011000101100 : romData <= 32'h0100739E;
      12'b011000101101 : romData <= 32'hDAFFFF03;
      12'b011000101110 : romData <= 32'h0400319E;
      12'b011000101111 : romData <= 32'h00F0801B;
      12'b011000110000 : romData <= 32'h00F0401B;
      12'b011000110001 : romData <= 32'h78099C9F;
      12'b011000110010 : romData <= 32'hD00A5A9F;
      12'b011000110011 : romData <= 32'h00F0A018;
      12'b011000110100 : romData <= 32'hF721A59C;
      12'b011000110101 : romData <= 32'h04E09CE0;
      12'b011000110110 : romData <= 32'hA5FBFF07;
      12'b011000110111 : romData <= 32'h04D07AE0;
      12'b011000111000 : romData <= 32'h00F0A018;
      12'b011000111001 : romData <= 32'h0004201A;
      12'b011000111010 : romData <= 32'h00FCE01A;
      12'b011000111011 : romData <= 32'hA121A59C;
      12'b011000111100 : romData <= 32'h0005A01A;
      12'b011000111101 : romData <= 32'hFFFF20AF;
      12'b011000111110 : romData <= 32'h00007186;
      12'b011000111111 : romData <= 32'h00C813E4;
      12'b011001000000 : romData <= 32'h11000010;
      12'b011001000001 : romData <= 32'h00B871E2;
      12'b011001000010 : romData <= 32'h009801D4;
      12'b011001000011 : romData <= 32'h04E09CE0;
      12'b011001000100 : romData <= 32'h04D07AE0;
      12'b011001000101 : romData <= 32'h20A801D4;
      12'b011001000110 : romData <= 32'h1CB801D4;
      12'b011001000111 : romData <= 32'h188801D4;
      12'b011001001000 : romData <= 32'h0C2801D4;
      12'b011001001001 : romData <= 32'h92FBFF07;
      12'b011001001010 : romData <= 32'h109801D4;
      12'b011001001011 : romData <= 32'h97FAFF07;
      12'b011001001100 : romData <= 32'h10006184;
      12'b011001001101 : romData <= 32'h2000A186;
      12'b011001001110 : romData <= 32'h1C00E186;
      12'b011001001111 : romData <= 32'h18002186;
      12'b011001010000 : romData <= 32'h0C00A184;
      12'b011001010001 : romData <= 32'h0400319E;
      12'b011001010010 : romData <= 32'h00A831E4;
      12'b011001010011 : romData <= 32'hEBFFFF13;
      12'b011001010100 : romData <= 32'hFFFF20AF;
      12'b011001010101 : romData <= 32'h00F0A018;
      12'b011001010110 : romData <= 32'h90FFFF03;
      12'b011001010111 : romData <= 32'h1522A59C;
      12'b011001011000 : romData <= 32'h00F0001B;
      12'b011001011001 : romData <= 32'h00F0401B;
      12'b011001011010 : romData <= 32'hD00A389E;
      12'b011001011011 : romData <= 32'h78095A9F;
      12'b011001011100 : romData <= 32'h00F0A018;
      12'b011001011101 : romData <= 32'h048871E0;
      12'b011001011110 : romData <= 32'h3022A59C;
      12'b011001011111 : romData <= 32'h04D09AE0;
      12'b011001100000 : romData <= 32'h7BFBFF07;
      12'b011001100001 : romData <= 32'h0C8801D4;
      12'b011001100010 : romData <= 32'h00F0201A;
      12'b011001100011 : romData <= 32'h5222319E;
      12'b011001100100 : romData <= 32'h0000001B;
      12'b011001100101 : romData <= 32'h108801D4;
      12'b011001100110 : romData <= 32'h04D09AE0;
      12'b011001100111 : romData <= 32'h1000A184;
      12'b011001101000 : romData <= 32'h73FBFF07;
      12'b011001101001 : romData <= 32'h0C006184;
      12'b011001101010 : romData <= 32'h0000201A;
      12'b011001101011 : romData <= 32'h0002601A;
      12'b011001101100 : romData <= 32'h0200A0AA;
      12'b011001101101 : romData <= 32'h00A818E4;
      12'b011001101110 : romData <= 32'h03000010;
      12'b011001101111 : romData <= 32'h00000015;
      12'b011001110000 : romData <= 32'h0100F172;
      12'b011001110001 : romData <= 32'h008811D4;
      12'b011001110010 : romData <= 32'h0400319E;
      12'b011001110011 : romData <= 32'h009831E4;
      12'b011001110100 : romData <= 32'hF9FFFF13;
      12'b011001110101 : romData <= 32'h0200A0AA;
      12'b011001110110 : romData <= 32'h00F0A018;
      12'b011001110111 : romData <= 32'h5E22A59C;
      12'b011001111000 : romData <= 32'h04D09AE0;
      12'b011001111001 : romData <= 32'h62FBFF07;
      12'b011001111010 : romData <= 32'h0C006184;
      12'b011001111011 : romData <= 32'h0000201A;
      12'b011001111100 : romData <= 32'h0000801B;
      12'b011001111101 : romData <= 32'h0002E01A;
      12'b011001111110 : romData <= 32'h020060AA;
      12'b011001111111 : romData <= 32'h009818E4;
      12'b011010000000 : romData <= 32'h03000010;
      12'b011010000001 : romData <= 32'h00000015;
      12'b011010000010 : romData <= 32'h01003173;
      12'b011010000011 : romData <= 32'h00003187;
      12'b011010000100 : romData <= 32'h008819E4;
      12'b011010000101 : romData <= 32'h14000010;
      12'b011010000110 : romData <= 32'h1D0060AA;
      12'b011010000111 : romData <= 32'h00985CE4;
      12'b011010001000 : romData <= 32'h10000010;
      12'b011010001001 : romData <= 32'h01003C9F;
      12'b011010001010 : romData <= 32'h00007186;
      12'b011010001011 : romData <= 32'h04D09AE0;
      12'b011010001100 : romData <= 32'h088801D4;
      12'b011010001101 : romData <= 32'h008801D4;
      12'b011010001110 : romData <= 32'h049801D4;
      12'b011010001111 : romData <= 32'h20B801D4;
      12'b011010010000 : romData <= 32'h1CC801D4;
      12'b011010010001 : romData <= 32'h188801D4;
      12'b011010010010 : romData <= 32'h1400A184;
      12'b011010010011 : romData <= 32'h48FBFF07;
      12'b011010010100 : romData <= 32'h0C006184;
      12'b011010010101 : romData <= 32'h2000E186;
      12'b011010010110 : romData <= 32'h1C002187;
      12'b011010010111 : romData <= 32'h18002186;
      12'b011010011000 : romData <= 32'h04C899E3;
      12'b011010011001 : romData <= 32'h0400319E;
      12'b011010011010 : romData <= 32'h00B831E4;
      12'b011010011011 : romData <= 32'hE4FFFF13;
      12'b011010011100 : romData <= 32'h020060AA;
      12'b011010011101 : romData <= 32'h0000201A;
      12'b011010011110 : romData <= 32'h00881CE4;
      12'b011010011111 : romData <= 32'h11000010;
      12'b011010100000 : romData <= 32'h0100189F;
      12'b011010100001 : romData <= 32'hFFFF189F;
      12'b011010100010 : romData <= 32'h00F0A018;
      12'b011010100011 : romData <= 32'h00E001D4;
      12'b011010100100 : romData <= 32'h8822A59C;
      12'b011010100101 : romData <= 32'h04D09AE0;
      12'b011010100110 : romData <= 32'h35FBFF07;
      12'b011010100111 : romData <= 32'h0C006184;
      12'b011010101000 : romData <= 32'h00F0A018;
      12'b011010101001 : romData <= 32'h00E001D4;
      12'b011010101010 : romData <= 32'hA122A59C;
      12'b011010101011 : romData <= 32'h04D09AE0;
      12'b011010101100 : romData <= 32'h2FFBFF07;
      12'b011010101101 : romData <= 32'h0C006184;
      12'b011010101110 : romData <= 32'h76FDFF03;
      12'b011010101111 : romData <= 32'h0000001B;
      12'b011010110000 : romData <= 32'h030020AA;
      12'b011010110001 : romData <= 32'h008838E4;
      12'b011010110010 : romData <= 32'hB5FFFF13;
      12'b011010110011 : romData <= 32'h04D09AE0;
      12'b011010110100 : romData <= 32'hF5FFFF03;
      12'b011010110101 : romData <= 32'h00F0A018;
      12'b011010110110 : romData <= 32'h7F00401B;
      12'b011010110111 : romData <= 32'hFCFF5AAB;
      12'b011010111000 : romData <= 32'h00F08018;
      12'b011010111001 : romData <= 32'h00F06018;
      12'b011010111010 : romData <= 32'h00D02EE4;
      12'b011010111011 : romData <= 32'h7809849C;
      12'b011010111100 : romData <= 32'h08000010;
      12'b011010111101 : romData <= 32'hD00A639C;
      12'b011010111110 : romData <= 32'h00F0A018;
      12'b011010111111 : romData <= 32'hBC22A59C;
      12'b011011000000 : romData <= 32'h1BFBFF07;
      12'b011011000001 : romData <= 32'h00C0C019;
      12'b011011000010 : romData <= 32'h62FDFF03;
      12'b011011000011 : romData <= 32'hFC1FCEA9;
      12'b011011000100 : romData <= 32'h00F0A018;
      12'b011011000101 : romData <= 32'h16FBFF07;
      12'b011011000110 : romData <= 32'hD222A59C;
      12'b011011000111 : romData <= 32'h5DFDFF03;
      12'b011011001000 : romData <= 32'h04D0DAE1;
      12'b011011001001 : romData <= 32'hA3FBFF07;
      12'b011011001010 : romData <= 32'h00000015;
      12'b011011001011 : romData <= 32'hA1FBFF07;
      12'b011011001100 : romData <= 32'hFF004BA7;
      12'b011011001101 : romData <= 32'hD0FF5A9F;
      12'b011011001110 : romData <= 32'h020020AA;
      12'b011011001111 : romData <= 32'h08883AE2;
      12'b011011010000 : romData <= 32'hFF004BA6;
      12'b011011010001 : romData <= 32'h00D031E2;
      12'b011011010010 : romData <= 32'h008831E2;
      12'b011011010011 : romData <= 32'hD0FF529E;
      12'b011011010100 : romData <= 32'h50FDFF03;
      12'b011011010101 : romData <= 32'h008852E2;
      12'b011011010110 : romData <= 32'h01009C9F;
      12'b011011010111 : romData <= 32'h000160AA;
      12'b011011011000 : romData <= 32'h00983CE4;
      12'b011011011001 : romData <= 32'hB0FDFF13;
      12'b011011011010 : romData <= 32'h0300B59E;
      12'b011011011011 : romData <= 32'h00F0A018;
      12'b011011011100 : romData <= 32'h7823A59C;
      12'b011011011101 : romData <= 32'hDDFDFF03;
      12'b011011011110 : romData <= 32'h00008018;
      12'b011011011111 : romData <= 32'h00881EE4;
      12'b011011100000 : romData <= 32'h17000010;
      12'b011011100001 : romData <= 32'h080020AA;
      12'b011011100010 : romData <= 32'h0888D6E2;
      12'b011011100011 : romData <= 32'h0100DE9F;
      12'b011011100100 : romData <= 32'h040020AA;
      12'b011011100101 : romData <= 32'h00883EE4;
      12'b011011100110 : romData <= 32'h40000010;
      12'b011011100111 : romData <= 32'h00B0DCE2;
      12'b011011101000 : romData <= 32'h00D030E4;
      12'b011011101001 : romData <= 32'h10000010;
      12'b011011101010 : romData <= 32'hFF0F20AA;
      12'b011011101011 : romData <= 32'h008834E4;
      12'b011011101100 : romData <= 32'h4A000010;
      12'b011011101101 : romData <= 32'h00F0A018;
      12'b011011101110 : romData <= 32'h00F08018;
      12'b011011101111 : romData <= 32'h00F06018;
      12'b011011110000 : romData <= 32'hEA22A59C;
      12'b011011110001 : romData <= 32'h7809849C;
      12'b011011110010 : romData <= 32'hE9FAFF07;
      12'b011011110011 : romData <= 32'hD00A639C;
      12'b011011110100 : romData <= 32'h010040AA;
      12'b011011110101 : romData <= 32'h45000000;
      12'b011011110110 : romData <= 32'h001080AA;
      12'b011011110111 : romData <= 32'hECFFFF03;
      12'b011011111000 : romData <= 32'h0000C01A;
      12'b011011111001 : romData <= 32'h0004201A;
      12'b011011111010 : romData <= 32'h008830E4;
      12'b011011111011 : romData <= 32'h0E000010;
      12'b011011111100 : romData <= 32'h0000201A;
      12'b011011111101 : romData <= 32'h008834E4;
      12'b011011111110 : romData <= 32'h26FDFF13;
      12'b011011111111 : romData <= 32'h010040AA;
      12'b011100000000 : romData <= 32'h00F0A018;
      12'b011100000001 : romData <= 32'h00F08018;
      12'b011100000010 : romData <= 32'h00F06018;
      12'b011100000011 : romData <= 32'h1923A59C;
      12'b011100000100 : romData <= 32'h7809849C;
      12'b011100000101 : romData <= 32'hD6FAFF07;
      12'b011100000110 : romData <= 32'hD00A639C;
      12'b011100000111 : romData <= 32'h1DFDFF03;
      12'b011100001000 : romData <= 32'h049092E2;
      12'b011100001001 : romData <= 32'h020020AA;
      12'b011100001010 : romData <= 32'h0888D4E3;
      12'b011100001011 : romData <= 32'h0000601A;
      12'b011100001100 : romData <= 32'hFF3F34A6;
      12'b011100001101 : romData <= 32'h009831E4;
      12'b011100001110 : romData <= 32'h08000010;
      12'b011100001111 : romData <= 32'h00F0A018;
      12'b011100010000 : romData <= 32'h00F06018;
      12'b011100010001 : romData <= 32'h00F001D4;
      12'b011100010010 : romData <= 32'h3A23A59C;
      12'b011100010011 : romData <= 32'h00008018;
      12'b011100010100 : romData <= 32'hC7FAFF07;
      12'b011100010101 : romData <= 32'hD00A639C;
      12'b011100010110 : romData <= 32'h0000201A;
      12'b011100010111 : romData <= 32'h008802E4;
      12'b011100011000 : romData <= 32'h10000010;
      12'b011100011001 : romData <= 32'h00F030E2;
      12'b011100011010 : romData <= 32'h0100B672;
      12'b011100011011 : romData <= 32'h00A811D4;
      12'b011100011100 : romData <= 32'h0100949E;
      12'b011100011101 : romData <= 32'h00A078E4;
      12'b011100011110 : romData <= 32'h07000010;
      12'b011100011111 : romData <= 32'h0000201A;
      12'b011100100000 : romData <= 32'h008802E4;
      12'b011100100001 : romData <= 32'h03000010;
      12'b011100100010 : romData <= 32'h00000015;
      12'b011100100011 : romData <= 32'h04A010D4;
      12'b011100100100 : romData <= 32'h04A014E3;
      12'b011100100101 : romData <= 32'h0000C01B;
      12'b011100100110 : romData <= 32'h6FFDFF03;
      12'b011100100111 : romData <= 32'hFFFF529E;
      12'b011100101000 : romData <= 32'h00003186;
      12'b011100101001 : romData <= 32'h01003172;
      12'b011100101010 : romData <= 32'h008816E4;
      12'b011100101011 : romData <= 32'hF1FFFF13;
      12'b011100101100 : romData <= 32'h00008018;
      12'b011100101101 : romData <= 32'h00F06018;
      12'b011100101110 : romData <= 32'h08B001D4;
      12'b011100101111 : romData <= 32'h048801D4;
      12'b011100110000 : romData <= 32'h00F001D4;
      12'b011100110001 : romData <= 32'hD00A639C;
      12'b011100110010 : romData <= 32'hA9FAFF07;
      12'b011100110011 : romData <= 32'h0C00A184;
      12'b011100110100 : romData <= 32'hE9FFFF03;
      12'b011100110101 : romData <= 32'h0100949E;
      12'b011100110110 : romData <= 32'h008854E4;
      12'b011100110111 : romData <= 32'hD2FFFF0F;
      12'b011100111000 : romData <= 32'h00000015;
      12'b011100111001 : romData <= 32'h010040AA;
      12'b011100111010 : romData <= 32'hEAFCFF03;
      12'b011100111011 : romData <= 32'h0000001B;
      12'b011100111100 : romData <= 32'h20737562;
      12'b011100111101 : romData <= 32'h6F727265;
      12'b011100111110 : romData <= 32'h000A2172;
      12'b011100111111 : romData <= 32'h61746144;
      12'b011101000000 : romData <= 32'h67617020;
      12'b011101000001 : romData <= 32'h61662065;
      12'b011101000010 : romData <= 32'h0A746C75;
      12'b011101000011 : romData <= 32'h70206900;
      12'b011101000100 : romData <= 32'h20656761;
      12'b011101000101 : romData <= 32'h6C756166;
      12'b011101000110 : romData <= 32'h74000A74;
      12'b011101000111 : romData <= 32'h0A6B6369;
      12'b011101001000 : romData <= 32'h6C6C6100;
      12'b011101001001 : romData <= 32'h216E6769;
      12'b011101001010 : romData <= 32'h3F3F000A;
      12'b011101001011 : romData <= 32'h000A3F3F;
      12'b011101001100 : romData <= 32'h676E6970;
      12'b011101001101 : romData <= 32'h7464000A;
      12'b011101001110 : romData <= 32'h000A626C;
      12'b011101001111 : romData <= 32'h626C7469;
      12'b011101010000 : romData <= 32'h6152000A;
      12'b011101010001 : romData <= 32'h2165676E;
      12'b011101010010 : romData <= 32'h7953000A;
      12'b011101010011 : romData <= 32'h6C616373;
      12'b011101010100 : romData <= 32'h54000A6C;
      12'b011101010101 : romData <= 32'h21706172;
      12'b011101010110 : romData <= 32'h7242000A;
      12'b011101010111 : romData <= 32'h0A6B6165;
      12'b011101011000 : romData <= 32'h65684300;
      12'b011101011001 : romData <= 32'h6E696B63;
      12'b011101011010 : romData <= 32'h616C2067;
      12'b011101011011 : romData <= 32'h70207473;
      12'b011101011100 : romData <= 32'h20656761;
      12'b011101011101 : romData <= 32'h6620666F;
      12'b011101011110 : romData <= 32'h6873616C;
      12'b011101011111 : romData <= 32'h706D6520;
      12'b011101100000 : romData <= 32'h000A7974;
      12'b011101100001 : romData <= 32'h73616C46;
      12'b011101100010 : romData <= 32'h72652068;
      12'b011101100011 : romData <= 32'h21726F72;
      12'b011101100100 : romData <= 32'h7245000A;
      12'b011101100101 : romData <= 32'h6E697361;
      12'b011101100110 : romData <= 32'h616C2067;
      12'b011101100111 : romData <= 32'h70207473;
      12'b011101101000 : romData <= 32'h20656761;
      12'b011101101001 : romData <= 32'h4620666F;
      12'b011101101010 : romData <= 32'h6873616C;
      12'b011101101011 : romData <= 32'h7257000A;
      12'b011101101100 : romData <= 32'h6E697469;
      12'b011101101101 : romData <= 32'h65742067;
      12'b011101101110 : romData <= 32'h73207473;
      12'b011101101111 : romData <= 32'h65757165;
      12'b011101110000 : romData <= 32'h2065636E;
      12'b011101110001 : romData <= 32'h66206F74;
      12'b011101110010 : romData <= 32'h6873616C;
      12'b011101110011 : romData <= 32'h56000A2E;
      12'b011101110100 : romData <= 32'h66697265;
      12'b011101110101 : romData <= 32'h676E6979;
      12'b011101110110 : romData <= 32'h73657420;
      12'b011101110111 : romData <= 32'h65732074;
      12'b011101111000 : romData <= 32'h6E657571;
      12'b011101111001 : romData <= 32'h66206563;
      12'b011101111010 : romData <= 32'h206D6F72;
      12'b011101111011 : romData <= 32'h73616C66;
      12'b011101111100 : romData <= 32'h000A2E68;
      12'b011101111101 : romData <= 32'h74736554;
      12'b011101111110 : romData <= 32'h69616620;
      12'b011101111111 : romData <= 32'h3A64656C;
      12'b011110000000 : romData <= 32'h20642520;
      12'b011110000001 : romData <= 32'h7830203A;
      12'b011110000010 : romData <= 32'h2F205825;
      12'b011110000011 : romData <= 32'h7830203D;
      12'b011110000100 : romData <= 32'h000A5825;
      12'b011110000101 : romData <= 32'h73616C46;
      12'b011110000110 : romData <= 32'h65742068;
      12'b011110000111 : romData <= 32'h6F207473;
      12'b011110001000 : romData <= 32'h2E79616B;
      12'b011110001001 : romData <= 32'h53000A0A;
      12'b011110001010 : romData <= 32'h6D617264;
      12'b011110001011 : romData <= 32'h746F6E20;
      12'b011110001100 : romData <= 32'h726F7720;
      12'b011110001101 : romData <= 32'h676E696B;
      12'b011110001110 : romData <= 32'h726F6320;
      12'b011110001111 : romData <= 32'h74636572;
      12'b011110010000 : romData <= 32'h202C796C;
      12'b011110010001 : romData <= 32'h61656C70;
      12'b011110010010 : romData <= 32'h63206573;
      12'b011110010011 : romData <= 32'h676E6168;
      12'b011110010100 : romData <= 32'h6F792065;
      12'b011110010101 : romData <= 32'h62207275;
      12'b011110010110 : romData <= 32'h6472616F;
      12'b011110010111 : romData <= 32'h4A000A21;
      12'b011110011000 : romData <= 32'h69706D75;
      12'b011110011001 : romData <= 32'h7420676E;
      12'b011110011010 : romData <= 32'h7270206F;
      12'b011110011011 : romData <= 32'h6172676F;
      12'b011110011100 : romData <= 32'h40206D6D;
      12'b011110011101 : romData <= 32'h58257830;
      12'b011110011110 : romData <= 32'h5343000A;
      12'b011110011111 : romData <= 32'h3337342D;
      12'b011110100000 : romData <= 32'h73795320;
      12'b011110100001 : romData <= 32'h206D6574;
      12'b011110100010 : romData <= 32'h676F7270;
      12'b011110100011 : romData <= 32'h6D6D6172;
      12'b011110100100 : romData <= 32'h20676E69;
      12'b011110100101 : romData <= 32'h20726F66;
      12'b011110100110 : romData <= 32'h74737973;
      12'b011110100111 : romData <= 32'h20736D65;
      12'b011110101000 : romData <= 32'h63206E6F;
      12'b011110101001 : romData <= 32'h0A706968;
      12'b011110101010 : romData <= 32'h65704F00;
      12'b011110101011 : romData <= 32'h7369726E;
      12'b011110101100 : romData <= 32'h61622063;
      12'b011110101101 : romData <= 32'h20646573;
      12'b011110101110 : romData <= 32'h74726976;
      12'b011110101111 : romData <= 32'h206C6175;
      12'b011110110000 : romData <= 32'h746F7250;
      12'b011110110001 : romData <= 32'h7079746F;
      12'b011110110010 : romData <= 32'h000A2E65;
      12'b011110110011 : romData <= 32'h6C697542;
      12'b011110110100 : romData <= 32'h65762064;
      12'b011110110101 : romData <= 32'h6F697372;
      12'b011110110110 : romData <= 32'h53203A6E;
      12'b011110110111 : romData <= 32'h4A206E75;
      12'b011110111000 : romData <= 32'h32206C75;
      12'b011110111001 : romData <= 32'h30312037;
      12'b011110111010 : romData <= 32'h3A39313A;
      12'b011110111011 : romData <= 32'h41203534;
      12'b011110111100 : romData <= 32'h4543204D;
      12'b011110111101 : romData <= 32'h32205453;
      12'b011110111110 : romData <= 32'h0A353230;
      12'b011110111111 : romData <= 32'h2049000A;
      12'b011111000000 : romData <= 32'h43206D61;
      12'b011111000001 : romData <= 32'h25205550;
      12'b011111000010 : romData <= 32'h666F2064;
      12'b011111000011 : romData <= 32'h20642520;
      12'b011111000100 : romData <= 32'h6E6E7572;
      12'b011111000101 : romData <= 32'h20676E69;
      12'b011111000110 : romData <= 32'h00207461;
      12'b011111000111 : romData <= 32'h64256425;
      12'b011111001000 : romData <= 32'h2564252E;
      12'b011111001001 : romData <= 32'h484D2064;
      12'b011111001010 : romData <= 32'h0A0A2E7A;
      12'b011111001011 : romData <= 32'h69615700;
      12'b011111001100 : romData <= 32'h676E6974;
      12'b011111001101 : romData <= 32'h726F6620;
      12'b011111001110 : romData <= 32'h55504320;
      12'b011111001111 : romData <= 32'h74203120;
      12'b011111010000 : romData <= 32'h6361206F;
      12'b011111010001 : romData <= 32'h61766974;
      12'b011111010010 : romData <= 32'h6D206574;
      12'b011111010011 : romData <= 32'h4A000A65;
      12'b011111010100 : romData <= 32'h69706D75;
      12'b011111010101 : romData <= 32'h7420676E;
      12'b011111010110 : romData <= 32'h616D206F;
      12'b011111010111 : romData <= 32'h70206E69;
      12'b011111011000 : romData <= 32'h72676F72;
      12'b011111011001 : romData <= 32'h40206D61;
      12'b011111011010 : romData <= 32'h58257830;
      12'b011111011011 : romData <= 32'h7250000A;
      12'b011111011100 : romData <= 32'h6172676F;
      12'b011111011101 : romData <= 32'h7270206D;
      12'b011111011110 : romData <= 32'h6E657365;
      12'b011111011111 : romData <= 32'h75622074;
      12'b011111100000 : romData <= 32'h6F6E2074;
      12'b011111100001 : romData <= 32'h6F662074;
      12'b011111100010 : romData <= 32'h68742072;
      12'b011111100011 : romData <= 32'h54207369;
      12'b011111100100 : romData <= 32'h65677261;
      12'b011111100101 : romData <= 32'h440A2E74;
      12'b011111100110 : romData <= 32'h79206469;
      12'b011111100111 : romData <= 32'h7520756F;
      12'b011111101000 : romData <= 32'h616F6C70;
      12'b011111101001 : romData <= 32'h6F662064;
      12'b011111101010 : romData <= 32'h68742072;
      12'b011111101011 : romData <= 32'h524F2065;
      12'b011111101100 : romData <= 32'h30303331;
      12'b011111101101 : romData <= 32'h616C7020;
      12'b011111101110 : romData <= 32'h726F6674;
      12'b011111101111 : romData <= 32'h000A3F6D;
      12'b011111110000 : romData <= 32'h6E776F44;
      12'b011111110001 : romData <= 32'h64616F6C;
      12'b011111110010 : romData <= 32'h6F64203A;
      12'b011111110011 : romData <= 32'h000A656E;
      12'b011111110100 : romData <= 32'h64616552;
      12'b011111110101 : romData <= 32'h20676E69;
      12'b011111110110 : romData <= 32'h65646F63;
      12'b011111110111 : romData <= 32'h62617420;
      12'b011111111000 : romData <= 32'h000A656C;
      12'b011111111001 : romData <= 32'h6E776F44;
      12'b011111111010 : romData <= 32'h64616F6C;
      12'b011111111011 : romData <= 32'h6573203A;
      12'b011111111100 : romData <= 32'h64612074;
      12'b011111111101 : romData <= 32'h73657264;
      12'b011111111110 : romData <= 32'h203D2073;
      12'b011111111111 : romData <= 32'h58257830;
      12'b100000000000 : romData <= 32'h7245000A;
      12'b100000000001 : romData <= 32'h2C726F72;
      12'b100000000010 : romData <= 32'h206F6E20;
      12'b100000000011 : romData <= 32'h676F7270;
      12'b100000000100 : romData <= 32'h206D6172;
      12'b100000000101 : romData <= 32'h64616F6C;
      12'b100000000110 : romData <= 32'h0A216465;
      12'b100000000111 : romData <= 32'h6D754A00;
      12'b100000001000 : romData <= 32'h676E6970;
      12'b100000001001 : romData <= 32'h206F7420;
      12'b100000001010 : romData <= 32'h676F7270;
      12'b100000001011 : romData <= 32'h6D6D6172;
      12'b100000001100 : romData <= 32'h7245000A;
      12'b100000001101 : romData <= 32'h2C726F72;
      12'b100000001110 : romData <= 32'h206F6E20;
      12'b100000001111 : romData <= 32'h676F7270;
      12'b100000010000 : romData <= 32'h206D6172;
      12'b100000010001 : romData <= 32'h46206E69;
      12'b100000010010 : romData <= 32'h6873616C;
      12'b100000010011 : romData <= 32'h53000A21;
      12'b100000010100 : romData <= 32'h69747465;
      12'b100000010101 : romData <= 32'h7020676E;
      12'b100000010110 : romData <= 32'h2E676F72;
      12'b100000010111 : romData <= 32'h646F6D20;
      12'b100000011000 : romData <= 32'h53000A65;
      12'b100000011001 : romData <= 32'h69747465;
      12'b100000011010 : romData <= 32'h7620676E;
      12'b100000011011 : romData <= 32'h66697265;
      12'b100000011100 : romData <= 32'h6F6D202E;
      12'b100000011101 : romData <= 32'h000A6564;
      12'b100000011110 : romData <= 32'h70206F4E;
      12'b100000011111 : romData <= 32'h72676F72;
      12'b100000100000 : romData <= 32'h70206D61;
      12'b100000100001 : romData <= 32'h65736572;
      12'b100000100010 : romData <= 32'h000A746E;
      12'b100000100011 : romData <= 32'h676F7250;
      12'b100000100100 : romData <= 32'h206D6172;
      12'b100000100101 : romData <= 32'h6D206E69;
      12'b100000100110 : romData <= 32'h66206D65;
      12'b100000100111 : romData <= 32'h206D6F72;
      12'b100000101000 : romData <= 32'h58257830;
      12'b100000101001 : romData <= 32'h206F7420;
      12'b100000101010 : romData <= 32'h58257830;
      12'b100000101011 : romData <= 32'h7753000A;
      12'b100000101100 : romData <= 32'h68637469;
      12'b100000101101 : romData <= 32'h74206465;
      12'b100000101110 : romData <= 32'h6F73206F;
      12'b100000101111 : romData <= 32'h622D7466;
      12'b100000110000 : romData <= 32'h0A736F69;
      12'b100000110001 : romData <= 32'h69775300;
      12'b100000110010 : romData <= 32'h65686374;
      12'b100000110011 : romData <= 32'h6F742064;
      12'b100000110100 : romData <= 32'h616C4620;
      12'b100000110101 : romData <= 32'h000A6873;
      12'b100000110110 : romData <= 32'h74697753;
      12'b100000110111 : romData <= 32'h64656863;
      12'b100000111000 : romData <= 32'h206F7420;
      12'b100000111001 : romData <= 32'h61524453;
      12'b100000111010 : romData <= 32'h50000A6D;
      12'b100000111011 : romData <= 32'h7361656C;
      12'b100000111100 : romData <= 32'h68632065;
      12'b100000111101 : romData <= 32'h65676E61;
      12'b100000111110 : romData <= 32'h206F7420;
      12'b100000111111 : romData <= 32'h20656874;
      12'b100001000000 : romData <= 32'h41524453;
      12'b100001000001 : romData <= 32'h7962204D;
      12'b100001000010 : romData <= 32'h0A742A20;
      12'b100001000011 : romData <= 32'h206F4E00;
      12'b100001000100 : romData <= 32'h676F7270;
      12'b100001000101 : romData <= 32'h206D6172;
      12'b100001000110 : romData <= 32'h64616F6C;
      12'b100001000111 : romData <= 32'h69206465;
      12'b100001001000 : romData <= 32'h4453206E;
      12'b100001001001 : romData <= 32'h216D6152;
      12'b100001001010 : romData <= 32'h7250000A;
      12'b100001001011 : romData <= 32'h6172676F;
      12'b100001001100 : romData <= 32'h6F64206D;
      12'b100001001101 : romData <= 32'h6E207365;
      12'b100001001110 : romData <= 32'h6620746F;
      12'b100001001111 : romData <= 32'h69207469;
      12'b100001010000 : romData <= 32'h6C46206E;
      12'b100001010001 : romData <= 32'h21687361;
      12'b100001010010 : romData <= 32'h6F43000A;
      12'b100001010011 : romData <= 32'h7261706D;
      12'b100001010100 : romData <= 32'h72652065;
      12'b100001010101 : romData <= 32'h20726F72;
      12'b100001010110 : romData <= 32'h30207461;
      12'b100001010111 : romData <= 32'h20582578;
      12'b100001011000 : romData <= 32'h7830203A;
      12'b100001011001 : romData <= 32'h21205825;
      12'b100001011010 : romData <= 32'h7830203D;
      12'b100001011011 : romData <= 32'h000A5825;
      12'b100001011100 : romData <= 32'h706D6F43;
      12'b100001011101 : romData <= 32'h20657261;
      12'b100001011110 : romData <= 32'h656E6F64;
      12'b100001011111 : romData <= 32'h6843000A;
      12'b100001100000 : romData <= 32'h696B6365;
      12'b100001100001 : romData <= 32'h6920676E;
      12'b100001100010 : romData <= 32'h68742066;
      12'b100001100011 : romData <= 32'h6C662065;
      12'b100001100100 : romData <= 32'h20687361;
      12'b100001100101 : romData <= 32'h65207369;
      12'b100001100110 : romData <= 32'h7974706D;
      12'b100001100111 : romData <= 32'h0A2E2E2E;
      12'b100001101000 : romData <= 32'h61745300;
      12'b100001101001 : romData <= 32'h66207472;
      12'b100001101010 : romData <= 32'h6873616C;
      12'b100001101011 : romData <= 32'h61726520;
      12'b100001101100 : romData <= 32'h63206573;
      12'b100001101101 : romData <= 32'h656C6379;
      12'b100001101110 : romData <= 32'h726F6620;
      12'b100001101111 : romData <= 32'h67617020;
      12'b100001110000 : romData <= 32'h78302065;
      12'b100001110001 : romData <= 32'h000A5825;
      12'b100001110010 : romData <= 32'h72617453;
      12'b100001110011 : romData <= 32'h72702074;
      12'b100001110100 : romData <= 32'h6172676F;
      12'b100001110101 : romData <= 32'h6E696D6D;
      12'b100001110110 : romData <= 32'h6C662067;
      12'b100001110111 : romData <= 32'h0A687361;
      12'b100001111000 : romData <= 32'h6F725000;
      12'b100001111001 : romData <= 32'h6D617267;
      12'b100001111010 : romData <= 32'h676E696D;
      12'b100001111011 : romData <= 32'h6E696620;
      12'b100001111100 : romData <= 32'h65687369;
      12'b100001111101 : romData <= 32'h43000A64;
      12'b100001111110 : romData <= 32'h6B636568;
      12'b100001111111 : romData <= 32'h20676E69;
      12'b100010000000 : romData <= 32'h66206669;
      12'b100010000001 : romData <= 32'h6873616C;
      12'b100010000010 : romData <= 32'h20736920;
      12'b100010000011 : romData <= 32'h72696427;
      12'b100010000100 : romData <= 32'h0A277974;
      12'b100010000101 : romData <= 32'h616C4600;
      12'b100010000110 : romData <= 32'h69206873;
      12'b100010000111 : romData <= 32'h6D652073;
      12'b100010001000 : romData <= 32'h20797470;
      12'b100010001001 : romData <= 32'h61726528;
      12'b100010001010 : romData <= 32'h29646573;
      12'b100010001011 : romData <= 32'h000A0A2E;
      12'b100010001100 : romData <= 32'h72617453;
      12'b100010001101 : romData <= 32'h676E6974;
      12'b100010001110 : romData <= 32'h6D697320;
      12'b100010001111 : romData <= 32'h20656C70;
      12'b100010010000 : romData <= 32'h61524453;
      12'b100010010001 : romData <= 32'h656D206D;
      12'b100010010010 : romData <= 32'h6568636D;
      12'b100010010011 : romData <= 32'h0A2E6B63;
      12'b100010010100 : romData <= 32'h7257000A;
      12'b100010010101 : romData <= 32'h6E697469;
      12'b100010010110 : romData <= 32'h2E2E2E67;
      12'b100010010111 : romData <= 32'h6556000A;
      12'b100010011000 : romData <= 32'h79666972;
      12'b100010011001 : romData <= 32'h2E676E69;
      12'b100010011010 : romData <= 32'h000A2E2E;
      12'b100010011011 : romData <= 32'h6F727245;
      12'b100010011100 : romData <= 32'h30402072;
      12'b100010011101 : romData <= 32'h20582578;
      12'b100010011110 : romData <= 32'h7830203A;
      12'b100010011111 : romData <= 32'h21205825;
      12'b100010100000 : romData <= 32'h7830203D;
      12'b100010100001 : romData <= 32'h000A5825;
      12'b100010100010 : romData <= 32'h6F20724E;
      12'b100010100011 : romData <= 32'h72652066;
      12'b100010100100 : romData <= 32'h73726F72;
      12'b100010100101 : romData <= 32'h756F6620;
      12'b100010100110 : romData <= 32'h3A20646E;
      12'b100010100111 : romData <= 32'h0A642520;
      12'b100010101000 : romData <= 32'h6D654D00;
      12'b100010101001 : romData <= 32'h63656863;
      12'b100010101010 : romData <= 32'h6F64206B;
      12'b100010101011 : romData <= 32'h202C656E;
      12'b100010101100 : romData <= 32'h65206425;
      12'b100010101101 : romData <= 32'h726F7272;
      12'b100010101110 : romData <= 32'h000A0A73;
      12'b100010101111 : romData <= 32'h74746553;
      12'b100010110000 : romData <= 32'h20676E69;
      12'b100010110001 : romData <= 32'h63617473;
      12'b100010110010 : romData <= 32'h6F74206B;
      12'b100010110011 : romData <= 32'h4D505320;
      12'b100010110100 : romData <= 32'h6553000A;
      12'b100010110101 : romData <= 32'h6E697474;
      12'b100010110110 : romData <= 32'h74732067;
      12'b100010110111 : romData <= 32'h206B6361;
      12'b100010111000 : romData <= 32'h53206F74;
      12'b100010111001 : romData <= 32'h4D415244;
      12'b100010111010 : romData <= 32'h7250000A;
      12'b100010111011 : romData <= 32'h6172676F;
      12'b100010111100 : romData <= 32'h6F74206D;
      12'b100010111101 : romData <= 32'h6962206F;
      12'b100010111110 : romData <= 32'h6F742067;
      12'b100010111111 : romData <= 32'h74696620;
      12'b100011000000 : romData <= 32'h206E6920;
      12'b100011000001 : romData <= 32'h74666F53;
      12'b100011000010 : romData <= 32'h736F6962;
      12'b100011000011 : romData <= 32'h6261202C;
      12'b100011000100 : romData <= 32'h6974726F;
      12'b100011000101 : romData <= 32'h0A21676E;
      12'b100011000110 : romData <= 32'h6E614300;
      12'b100011000111 : romData <= 32'h20746F6E;
      12'b100011001000 : romData <= 32'h676F7270;
      12'b100011001001 : romData <= 32'h206D6172;
      12'b100011001010 : romData <= 32'h73616C66;
      12'b100011001011 : romData <= 32'h61202C68;
      12'b100011001100 : romData <= 32'h74726F62;
      12'b100011001101 : romData <= 32'h21676E69;
      12'b100011001110 : romData <= 32'h6F44000A;
      12'b100011001111 : romData <= 32'h6F6C6E77;
      12'b100011010000 : romData <= 32'h203A6461;
      12'b100011010001 : romData <= 32'h30207461;
      12'b100011010010 : romData <= 32'h0A582578;
      12'b100011010011 : romData <= 32'h72655600;
      12'b100011010100 : romData <= 32'h63696669;
      12'b100011010101 : romData <= 32'h6F697461;
      12'b100011010110 : romData <= 32'h7265206E;
      12'b100011010111 : romData <= 32'h20726F72;
      12'b100011011000 : romData <= 32'h30207461;
      12'b100011011001 : romData <= 32'h20582578;
      12'b100011011010 : romData <= 32'h7830203A;
      12'b100011011011 : romData <= 32'h21205825;
      12'b100011011100 : romData <= 32'h7830203D;
      12'b100011011101 : romData <= 32'h000A5825;
      12'b100011011110 : romData <= 32'h6E6B6E55;
      12'b100011011111 : romData <= 32'h206E776F;
      12'b100011100000 : romData <= 32'h65646F63;
      12'b100011100001 : romData <= 32'h6E4B0021;
      12'b100011100010 : romData <= 32'h206E776F;
      12'b100011100011 : romData <= 32'h33325352;
      12'b100011100100 : romData <= 32'h6F632032;
      12'b100011100101 : romData <= 32'h6E616D6D;
      12'b100011100110 : romData <= 32'h0A3A7364;
      12'b100011100111 : romData <= 32'h202A2A00;
      12'b100011101000 : romData <= 32'h72617453;
      12'b100011101001 : romData <= 32'h68742074;
      12'b100011101010 : romData <= 32'h72702065;
      12'b100011101011 : romData <= 32'h6172676F;
      12'b100011101100 : romData <= 32'h6F6C206D;
      12'b100011101101 : romData <= 32'h64656461;
      12'b100011101110 : romData <= 32'h206E6920;
      12'b100011101111 : romData <= 32'h67726174;
      12'b100011110000 : romData <= 32'h000A7465;
      12'b100011110001 : romData <= 32'h5320702A;
      12'b100011110010 : romData <= 32'h70207465;
      12'b100011110011 : romData <= 32'h72676F72;
      12'b100011110100 : romData <= 32'h696D6D61;
      12'b100011110101 : romData <= 32'h6D20676E;
      12'b100011110110 : romData <= 32'h2065646F;
      12'b100011110111 : romData <= 32'h66656428;
      12'b100011111000 : romData <= 32'h746C7561;
      12'b100011111001 : romData <= 32'h2A000A29;
      12'b100011111010 : romData <= 32'h65532076;
      12'b100011111011 : romData <= 32'h65762074;
      12'b100011111100 : romData <= 32'h69666972;
      12'b100011111101 : romData <= 32'h69746163;
      12'b100011111110 : romData <= 32'h6D206E6F;
      12'b100011111111 : romData <= 32'h0A65646F;
      12'b100100000000 : romData <= 32'h20692A00;
      12'b100100000001 : romData <= 32'h776F6853;
      12'b100100000010 : romData <= 32'h666E6920;
      12'b100100000011 : romData <= 32'h6E6F206F;
      12'b100100000100 : romData <= 32'h6F727020;
      12'b100100000101 : romData <= 32'h6D617267;
      12'b100100000110 : romData <= 32'h206E6920;
      12'b100100000111 : romData <= 32'h67726174;
      12'b100100001000 : romData <= 32'h000A7465;
      12'b100100001001 : romData <= 32'h5420742A;
      12'b100100001010 : romData <= 32'h6C67676F;
      12'b100100001011 : romData <= 32'h61742065;
      12'b100100001100 : romData <= 32'h74656772;
      12'b100100001101 : romData <= 32'h74656220;
      12'b100100001110 : romData <= 32'h6E656577;
      12'b100100001111 : romData <= 32'h52445320;
      12'b100100010000 : romData <= 32'h28206D61;
      12'b100100010001 : romData <= 32'h61666564;
      12'b100100010010 : romData <= 32'h29746C75;
      12'b100100010011 : romData <= 32'h6F73202C;
      12'b100100010100 : romData <= 32'h422D7466;
      12'b100100010101 : romData <= 32'h20736F69;
      12'b100100010110 : romData <= 32'h20646E61;
      12'b100100010111 : romData <= 32'h73616C46;
      12'b100100011000 : romData <= 32'h2A000A68;
      12'b100100011001 : romData <= 32'h6550206D;
      12'b100100011010 : romData <= 32'h726F6672;
      12'b100100011011 : romData <= 32'h6973206D;
      12'b100100011100 : romData <= 32'h656C706D;
      12'b100100011101 : romData <= 32'h52445320;
      12'b100100011110 : romData <= 32'h6D206D61;
      12'b100100011111 : romData <= 32'h68636D65;
      12'b100100100000 : romData <= 32'h0A6B6365;
      12'b100100100001 : romData <= 32'h20732A00;
      12'b100100100010 : romData <= 32'h63656843;
      12'b100100100011 : romData <= 32'h5053206B;
      12'b100100100100 : romData <= 32'h6C662D49;
      12'b100100100101 : romData <= 32'h20687361;
      12'b100100100110 : romData <= 32'h70696863;
      12'b100100100111 : romData <= 32'h652A000A;
      12'b100100101000 : romData <= 32'h61724520;
      12'b100100101001 : romData <= 32'h53206573;
      12'b100100101010 : romData <= 32'h462D4950;
      12'b100100101011 : romData <= 32'h6873616C;
      12'b100100101100 : romData <= 32'h69686320;
      12'b100100101101 : romData <= 32'h2A000A70;
      12'b100100101110 : romData <= 32'h74532066;
      12'b100100101111 : romData <= 32'h2065726F;
      12'b100100110000 : romData <= 32'h676F7270;
      12'b100100110001 : romData <= 32'h206D6172;
      12'b100100110010 : romData <= 32'h64616F6C;
      12'b100100110011 : romData <= 32'h69206465;
      12'b100100110100 : romData <= 32'h4453206E;
      12'b100100110101 : romData <= 32'h204D4152;
      12'b100100110110 : romData <= 32'h53206F74;
      12'b100100110111 : romData <= 32'h462D4950;
      12'b100100111000 : romData <= 32'h6873616C;
      12'b100100111001 : romData <= 32'h632A000A;
      12'b100100111010 : romData <= 32'h6D6F4320;
      12'b100100111011 : romData <= 32'h65726170;
      12'b100100111100 : romData <= 32'h6F727020;
      12'b100100111101 : romData <= 32'h6D617267;
      12'b100100111110 : romData <= 32'h616F6C20;
      12'b100100111111 : romData <= 32'h20646564;
      12'b100101000000 : romData <= 32'h53206E69;
      12'b100101000001 : romData <= 32'h4D415244;
      12'b100101000010 : romData <= 32'h74697720;
      12'b100101000011 : romData <= 32'h50532068;
      12'b100101000100 : romData <= 32'h6C462D49;
      12'b100101000101 : romData <= 32'h0A687361;
      12'b100101000110 : romData <= 32'h20722A00;
      12'b100101000111 : romData <= 32'h206E7552;
      12'b100101001000 : romData <= 32'h676F7270;
      12'b100101001001 : romData <= 32'h206D6172;
      12'b100101001010 : romData <= 32'h726F7473;
      12'b100101001011 : romData <= 32'h69206465;
      12'b100101001100 : romData <= 32'h5053206E;
      12'b100101001101 : romData <= 32'h6C462D49;
      12'b100101001110 : romData <= 32'h0A687361;
      12'b100101001111 : romData <= 32'h20712A00;
      12'b100101010000 : romData <= 32'h67676F54;
      12'b100101010001 : romData <= 32'h7320656C;
      12'b100101010010 : romData <= 32'h6B636174;
      12'b100101010011 : romData <= 32'h696F7020;
      12'b100101010100 : romData <= 32'h7265746E;
      12'b100101010101 : romData <= 32'h6F726620;
      12'b100101010110 : romData <= 32'h4453206D;
      12'b100101010111 : romData <= 32'h204D4152;
      12'b100101011000 : romData <= 32'h66656428;
      12'b100101011001 : romData <= 32'h746C7561;
      12'b100101011010 : romData <= 32'h69772029;
      12'b100101011011 : romData <= 32'h53206874;
      12'b100101011100 : romData <= 32'h000A4D50;
      12'b100101011101 : romData <= 32'h5420682A;
      12'b100101011110 : romData <= 32'h20736968;
      12'b100101011111 : romData <= 32'h706C6568;
      12'b100101100000 : romData <= 32'h65726373;
      12'b100101100001 : romData <= 32'h0A0A6E65;
      12'b100101100011 : romData <= 32'hEFBEADDE;
      12'b100101100100 : romData <= 32'h01000000;
      12'b100101100101 : romData <= 32'h02000000;
      12'b100101100110 : romData <= 32'h03000000;
      12'b100101100111 : romData <= 32'h04000000;
      12'b100101101000 : romData <= 32'h05000000;
      12'b100101101001 : romData <= 32'h06000000;
      12'b100101101010 : romData <= 32'h07000000;
      12'b100101101011 : romData <= 32'h862300F0;
      12'b100101101100 : romData <= 32'h9D2300F0;
      12'b100101101101 : romData <= 32'hC42300F0;
      12'b100101101110 : romData <= 32'hE72300F0;
      12'b100101101111 : romData <= 32'h012400F0;
      12'b100101110000 : romData <= 32'h242400F0;
      12'b100101110001 : romData <= 32'h632400F0;
      12'b100101110010 : romData <= 32'h852400F0;
      12'b100101110011 : romData <= 32'h9E2400F0;
      12'b100101110100 : romData <= 32'hB72400F0;
      12'b100101110101 : romData <= 32'hE62400F0;
      12'b100101110110 : romData <= 32'h192500F0;
      12'b100101110111 : romData <= 32'h3D2500F0;
      12'b100101111000 : romData <= 32'h742500F0;
      default : romData <= 32'd0;
    endcase

endmodule

